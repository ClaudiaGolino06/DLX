
library IEEE;

use IEEE.std_logic_1164.all;

package CONV_PACK_DLX_IR_SIZE32_PC_SIZE32 is

-- define attributes
attribute ENUM_ENCODING : STRING;

-- define any necessary types
type aluOp is (NOP, ADDS, LLS, LRS, ADD, SUB, ANDR, ORR, XORR, SNE, SLE, SGE, 
   BEQZ, BNEZ, SUBI, ANDI, ORI, XORI, SLLI, SRLI, SNEI, SLEI, SGEI, LW, SW, 
   SUBU, SUBUI, ADDU, ADDUI, SRA1, SEQ, SLT, SGT, SLTU, SGTU, SGEU, LHI, JR, 
   JALR, SRAI, SEQI, SLTI, SGTI, LB, LBU, LHU, SB, SLTUI, SGTUI, SGEUI, trap, 
   rfe);
attribute ENUM_ENCODING of aluOp : type is 
   "000000 000001 000010 000011 000100 000101 000110 000111 001000 001001 001010 001011 001100 001101 001110 001111 010000 010001 010010 010011 010100 010101 010110 010111 011000 011001 011010 011011 011100 011101 011110 011111 100000 100001 100010 100011 100100 100101 100110 100111 101000 101001 101010 101011 101100 101101 101110 101111 110000 110001 110010 110011";
   
   -- Declarations for conversion functions.
   function std_logic_vector_to_aluOp(arg : in std_logic_vector( 1 to 6 )) 
               return aluOp;
   function aluOp_to_std_logic_vector(arg : in aluOp) return std_logic_vector;

end CONV_PACK_DLX_IR_SIZE32_PC_SIZE32;

package body CONV_PACK_DLX_IR_SIZE32_PC_SIZE32 is
   
   -- std_logic_vector to enum type function
   function std_logic_vector_to_aluOp(arg : in std_logic_vector( 1 to 6 )) 
   return aluOp is
   -- synopsys built_in SYN_FEED_THRU;
   begin
      case arg is
         when "000000" => return NOP;
         when "000001" => return ADDS;
         when "000010" => return LLS;
         when "000011" => return LRS;
         when "000100" => return ADD;
         when "000101" => return SUB;
         when "000110" => return ANDR;
         when "000111" => return ORR;
         when "001000" => return XORR;
         when "001001" => return SNE;
         when "001010" => return SLE;
         when "001011" => return SGE;
         when "001100" => return BEQZ;
         when "001101" => return BNEZ;
         when "001110" => return SUBI;
         when "001111" => return ANDI;
         when "010000" => return ORI;
         when "010001" => return XORI;
         when "010010" => return SLLI;
         when "010011" => return SRLI;
         when "010100" => return SNEI;
         when "010101" => return SLEI;
         when "010110" => return SGEI;
         when "010111" => return LW;
         when "011000" => return SW;
         when "011001" => return SUBU;
         when "011010" => return SUBUI;
         when "011011" => return ADDU;
         when "011100" => return ADDUI;
         when "011101" => return SRA1;
         when "011110" => return SEQ;
         when "011111" => return SLT;
         when "100000" => return SGT;
         when "100001" => return SLTU;
         when "100010" => return SGTU;
         when "100011" => return SGEU;
         when "100100" => return LHI;
         when "100101" => return JR;
         when "100110" => return JALR;
         when "100111" => return SRAI;
         when "101000" => return SEQI;
         when "101001" => return SLTI;
         when "101010" => return SGTI;
         when "101011" => return LB;
         when "101100" => return LBU;
         when "101101" => return LHU;
         when "101110" => return SB;
         when "101111" => return SLTUI;
         when "110000" => return SGTUI;
         when "110001" => return SGEUI;
         when "110010" => return trap;
         when "110011" => return rfe;
         when others => assert FALSE -- this should not happen.
               report "un-convertible value"
               severity warning;
               return NOP;
      end case;
   end;
   
   -- enum type to std_logic_vector function
   function aluOp_to_std_logic_vector(arg : in aluOp) return std_logic_vector 
   is
   -- synopsys built_in SYN_FEED_THRU;
   begin
      case arg is
         when NOP => return "000000";
         when ADDS => return "000001";
         when LLS => return "000010";
         when LRS => return "000011";
         when ADD => return "000100";
         when SUB => return "000101";
         when ANDR => return "000110";
         when ORR => return "000111";
         when XORR => return "001000";
         when SNE => return "001001";
         when SLE => return "001010";
         when SGE => return "001011";
         when BEQZ => return "001100";
         when BNEZ => return "001101";
         when SUBI => return "001110";
         when ANDI => return "001111";
         when ORI => return "010000";
         when XORI => return "010001";
         when SLLI => return "010010";
         when SRLI => return "010011";
         when SNEI => return "010100";
         when SLEI => return "010101";
         when SGEI => return "010110";
         when LW => return "010111";
         when SW => return "011000";
         when SUBU => return "011001";
         when SUBUI => return "011010";
         when ADDU => return "011011";
         when ADDUI => return "011100";
         when SRA1 => return "011101";
         when SEQ => return "011110";
         when SLT => return "011111";
         when SGT => return "100000";
         when SLTU => return "100001";
         when SGTU => return "100010";
         when SGEU => return "100011";
         when LHI => return "100100";
         when JR => return "100101";
         when JALR => return "100110";
         when SRAI => return "100111";
         when SEQI => return "101000";
         when SLTI => return "101001";
         when SGTI => return "101010";
         when LB => return "101011";
         when LBU => return "101100";
         when LHU => return "101101";
         when SB => return "101110";
         when SLTUI => return "101111";
         when SGTUI => return "110000";
         when SGEUI => return "110001";
         when trap => return "110010";
         when rfe => return "110011";
         when others => assert FALSE -- this should not happen.
               report "un-convertible value"
               severity warning;
               return "000000";
      end case;
   end;

end CONV_PACK_DLX_IR_SIZE32_PC_SIZE32;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity 
   dlx_cu_MICROCODE_MEM_SIZE62_FUNC_SIZE11_OP_CODE_SIZE6_IR_SIZE32_CW_SIZE15_DW01_inc_5 
   is

   port( A : in std_logic_vector (31 downto 0);  SUM : out std_logic_vector (31
         downto 0));

end 
   dlx_cu_MICROCODE_MEM_SIZE62_FUNC_SIZE11_OP_CODE_SIZE6_IR_SIZE32_CW_SIZE15_DW01_inc_5;

architecture SYN_cla of 
   dlx_cu_MICROCODE_MEM_SIZE62_FUNC_SIZE11_OP_CODE_SIZE6_IR_SIZE32_CW_SIZE15_DW01_inc_5 
   is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      , n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, 
      n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45
      , n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, 
      n60, n61 : std_logic;

begin
   
   U2 : AND3_X1 port map( A1 => A(24), A2 => A(25), A3 => n9, ZN => n1);
   U3 : OR2_X1 port map( A1 => n43, A2 => n44, ZN => n2);
   U4 : NOR2_X1 port map( A1 => n52, A2 => n8, ZN => n7);
   U5 : NAND2_X1 port map( A1 => n3, A2 => n4, ZN => n40);
   U6 : AND2_X1 port map( A1 => n54, A2 => n55, ZN => n3);
   U7 : NOR2_X1 port map( A1 => n2, A2 => n8, ZN => n4);
   U8 : NOR2_X1 port map( A1 => n40, A2 => n10, ZN => n9);
   U9 : NOR2_X1 port map( A1 => n31, A2 => n32, ZN => n30);
   U10 : NOR2_X1 port map( A1 => n56, A2 => n57, ZN => n55);
   U11 : NAND2_X1 port map( A1 => n17, A2 => n59, ZN => n13);
   U12 : NOR2_X1 port map( A1 => n60, A2 => n61, ZN => n59);
   U13 : XNOR2_X1 port map( A => A(6), B => n16, ZN => SUM(6));
   U14 : XNOR2_X1 port map( A => A(14), B => n51, ZN => SUM(14));
   U15 : XNOR2_X1 port map( A => A(22), B => n39, ZN => SUM(22));
   U16 : XOR2_X1 port map( A => n6, B => A(10), Z => SUM(10));
   U17 : XOR2_X1 port map( A => n26, B => A(30), Z => SUM(30));
   U18 : XOR2_X1 port map( A => n5, B => A(18), Z => SUM(18));
   U19 : XOR2_X1 port map( A => n1, B => A(26), Z => SUM(26));
   U20 : XOR2_X1 port map( A => A(16), B => n7, Z => SUM(16));
   U21 : INV_X1 port map( A => n22, ZN => n21);
   U22 : XOR2_X1 port map( A => n23, B => A(31), Z => SUM(31));
   U23 : XOR2_X1 port map( A => n28, B => A(29), Z => SUM(29));
   U24 : XNOR2_X1 port map( A => A(5), B => n18, ZN => SUM(5));
   U25 : NAND2_X1 port map( A1 => A(4), A2 => n17, ZN => n18);
   U26 : XNOR2_X1 port map( A => A(9), B => n12, ZN => SUM(9));
   U27 : NAND2_X1 port map( A1 => A(8), A2 => n54, ZN => n12);
   U28 : XNOR2_X1 port map( A => A(13), B => n53, ZN => SUM(13));
   U29 : NAND2_X1 port map( A1 => A(12), A2 => n3, ZN => n53);
   U30 : XNOR2_X1 port map( A => A(17), B => n46, ZN => SUM(17));
   U31 : NAND2_X1 port map( A1 => A(16), A2 => n7, ZN => n46);
   U32 : XNOR2_X1 port map( A => A(21), B => n41, ZN => SUM(21));
   U33 : NAND2_X1 port map( A1 => A(20), A2 => n42, ZN => n41);
   U34 : XNOR2_X1 port map( A => A(25), B => n34, ZN => SUM(25));
   U35 : AND3_X1 port map( A1 => A(16), A2 => A(17), A3 => n7, ZN => n5);
   U36 : AND3_X1 port map( A1 => A(8), A2 => A(9), A3 => n54, ZN => n6);
   U37 : INV_X1 port map( A => A(28), ZN => n29);
   U38 : OR2_X1 port map( A1 => n47, A2 => n48, ZN => n8);
   U39 : NAND2_X1 port map( A1 => n54, A2 => n55, ZN => n52);
   U40 : XNOR2_X1 port map( A => A(3), B => n20, ZN => SUM(3));
   U41 : NAND2_X1 port map( A1 => A(24), A2 => n9, ZN => n34);
   U42 : INV_X1 port map( A => n9, ZN => n33);
   U43 : OR2_X1 port map( A1 => n35, A2 => n36, ZN => n10);
   U44 : XNOR2_X1 port map( A => A(20), B => n40, ZN => SUM(20));
   U45 : INV_X1 port map( A => n40, ZN => n42);
   U46 : XNOR2_X1 port map( A => A(12), B => n52, ZN => SUM(12));
   U47 : XOR2_X1 port map( A => A(27), B => n11, Z => SUM(27));
   U48 : AND2_X1 port map( A1 => n1, A2 => A(26), ZN => n11);
   U49 : XNOR2_X1 port map( A => A(8), B => n13, ZN => SUM(8));
   U50 : XNOR2_X1 port map( A => A(24), B => n33, ZN => SUM(24));
   U51 : NAND2_X1 port map( A1 => n9, A2 => n30, ZN => n25);
   U52 : XNOR2_X1 port map( A => A(2), B => n22, ZN => SUM(2));
   U53 : XNOR2_X1 port map( A => A(28), B => n25, ZN => SUM(28));
   U54 : NAND2_X1 port map( A1 => A(2), A2 => n21, ZN => n20);
   U55 : NOR2_X1 port map( A1 => n25, A2 => n29, ZN => n28);
   U56 : NOR2_X1 port map( A1 => n25, A2 => n27, ZN => n26);
   U57 : NOR2_X1 port map( A1 => n24, A2 => n25, ZN => n23);
   U58 : INV_X1 port map( A => A(0), ZN => SUM(0));
   U59 : NAND2_X1 port map( A1 => A(1), A2 => A(0), ZN => n22);
   U60 : NAND4_X1 port map( A1 => A(0), A2 => A(2), A3 => A(1), A4 => A(3), ZN 
                           => n19);
   U61 : XNOR2_X1 port map( A => A(7), B => n14, ZN => SUM(7));
   U62 : NAND2_X1 port map( A1 => n15, A2 => A(6), ZN => n14);
   U63 : INV_X1 port map( A => n16, ZN => n15);
   U64 : NAND3_X1 port map( A1 => A(4), A2 => A(5), A3 => n17, ZN => n16);
   U65 : XNOR2_X1 port map( A => A(4), B => n19, ZN => SUM(4));
   U66 : NAND3_X1 port map( A1 => A(30), A2 => A(29), A3 => A(28), ZN => n24);
   U67 : NAND2_X1 port map( A1 => A(28), A2 => A(29), ZN => n27);
   U68 : NAND2_X1 port map( A1 => A(24), A2 => A(25), ZN => n32);
   U69 : NAND2_X1 port map( A1 => A(27), A2 => A(26), ZN => n31);
   U70 : NAND2_X1 port map( A1 => A(20), A2 => A(21), ZN => n36);
   U71 : NAND2_X1 port map( A1 => A(23), A2 => A(22), ZN => n35);
   U72 : XNOR2_X1 port map( A => A(23), B => n37, ZN => SUM(23));
   U73 : NAND2_X1 port map( A1 => n38, A2 => A(22), ZN => n37);
   U74 : INV_X1 port map( A => n39, ZN => n38);
   U75 : NAND3_X1 port map( A1 => A(20), A2 => A(21), A3 => n42, ZN => n39);
   U76 : NAND2_X1 port map( A1 => A(16), A2 => A(17), ZN => n44);
   U77 : NAND2_X1 port map( A1 => A(19), A2 => A(18), ZN => n43);
   U78 : XOR2_X1 port map( A => A(1), B => A(0), Z => SUM(1));
   U79 : XNOR2_X1 port map( A => A(19), B => n45, ZN => SUM(19));
   U80 : NAND2_X1 port map( A1 => n5, A2 => A(18), ZN => n45);
   U81 : NAND2_X1 port map( A1 => A(12), A2 => A(13), ZN => n48);
   U82 : NAND2_X1 port map( A1 => A(15), A2 => A(14), ZN => n47);
   U83 : XNOR2_X1 port map( A => A(15), B => n49, ZN => SUM(15));
   U84 : NAND2_X1 port map( A1 => n50, A2 => A(14), ZN => n49);
   U85 : INV_X1 port map( A => n51, ZN => n50);
   U86 : NAND3_X1 port map( A1 => A(12), A2 => A(13), A3 => n3, ZN => n51);
   U87 : NAND2_X1 port map( A1 => A(8), A2 => A(9), ZN => n57);
   U88 : NAND2_X1 port map( A1 => A(11), A2 => A(10), ZN => n56);
   U89 : XNOR2_X1 port map( A => A(11), B => n58, ZN => SUM(11));
   U90 : NAND2_X1 port map( A1 => n6, A2 => A(10), ZN => n58);
   U91 : INV_X1 port map( A => n13, ZN => n54);
   U92 : NAND2_X1 port map( A1 => A(4), A2 => A(5), ZN => n61);
   U93 : NAND2_X1 port map( A1 => A(7), A2 => A(6), ZN => n60);
   U94 : INV_X1 port map( A => n19, ZN => n17);

end SYN_cla;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity 
   dlx_cu_MICROCODE_MEM_SIZE62_FUNC_SIZE11_OP_CODE_SIZE6_IR_SIZE32_CW_SIZE15_DW01_inc_4 
   is

   port( A : in std_logic_vector (31 downto 0);  SUM : out std_logic_vector (31
         downto 0));

end 
   dlx_cu_MICROCODE_MEM_SIZE62_FUNC_SIZE11_OP_CODE_SIZE6_IR_SIZE32_CW_SIZE15_DW01_inc_4;

architecture SYN_cla of 
   dlx_cu_MICROCODE_MEM_SIZE62_FUNC_SIZE11_OP_CODE_SIZE6_IR_SIZE32_CW_SIZE15_DW01_inc_4 
   is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal SUM_31_port, SUM_30_port, SUM_29_port, SUM_28_port, SUM_27_port, 
      SUM_26_port, SUM_25_port, SUM_24_port, SUM_23_port, SUM_22_port, 
      SUM_21_port, SUM_20_port, SUM_19_port, SUM_18_port, SUM_17_port, 
      SUM_16_port, SUM_15_port, SUM_14_port, SUM_13_port, SUM_12_port, 
      SUM_11_port, SUM_10_port, SUM_9_port, SUM_8_port, SUM_7_port, SUM_6_port,
      SUM_5_port, SUM_4_port, SUM_3_port, SUM_2_port, SUM_1_port, SUM_0_port, 
      n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, 
      n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31
      , n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, 
      n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60
      , n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, 
      n75 : std_logic;

begin
   SUM <= ( SUM_31_port, SUM_30_port, SUM_29_port, SUM_28_port, SUM_27_port, 
      SUM_26_port, SUM_25_port, SUM_24_port, SUM_23_port, SUM_22_port, 
      SUM_21_port, SUM_20_port, SUM_19_port, SUM_18_port, SUM_17_port, 
      SUM_16_port, SUM_15_port, SUM_14_port, SUM_13_port, SUM_12_port, 
      SUM_11_port, SUM_10_port, SUM_9_port, SUM_8_port, SUM_7_port, SUM_6_port,
      SUM_5_port, SUM_4_port, SUM_3_port, SUM_2_port, SUM_1_port, SUM_0_port );
   
   U2 : AND2_X1 port map( A1 => A(20), A2 => A(21), ZN => n1);
   U3 : BUF_X1 port map( A => n14, Z => n2);
   U4 : NAND2_X1 port map( A1 => n3, A2 => n4, ZN => n41);
   U5 : AND2_X1 port map( A1 => n25, A2 => n26, ZN => n3);
   U6 : NOR2_X1 port map( A1 => n46, A2 => n47, ZN => n4);
   U7 : XOR2_X1 port map( A => A(25), B => n5, Z => SUM_25_port);
   U8 : AND2_X1 port map( A1 => A(24), A2 => n3, ZN => n5);
   U9 : CLKBUF_X1 port map( A => A(2), Z => n6);
   U10 : INV_X1 port map( A => n2, ZN => n68);
   U11 : INV_X1 port map( A => n63, ZN => n7);
   U12 : AND2_X1 port map( A1 => n30, A2 => n8, ZN => n25);
   U13 : NOR2_X1 port map( A1 => n19, A2 => n7, ZN => n8);
   U14 : INV_X1 port map( A => n30, ZN => n9);
   U15 : CLKBUF_X1 port map( A => A(5), Z => n10);
   U16 : NOR2_X1 port map( A1 => n31, A2 => n19, ZN => n14);
   U17 : AND2_X1 port map( A1 => n25, A2 => n26, ZN => n11);
   U18 : XOR2_X1 port map( A => A(15), B => n12, Z => SUM_15_port);
   U19 : AND2_X1 port map( A1 => n66, A2 => A(14), ZN => n12);
   U20 : INV_X1 port map( A => SUM_0_port, ZN => n13);
   U21 : NOR2_X1 port map( A1 => n31, A2 => n19, ZN => n15);
   U22 : CLKBUF_X1 port map( A => A(4), Z => n16);
   U23 : AND2_X1 port map( A1 => n55, A2 => n1, ZN => n51);
   U24 : AND4_X1 port map( A1 => A(3), A2 => A(2), A3 => A(1), A4 => A(0), ZN 
                           => n17);
   U25 : AND4_X1 port map( A1 => A(1), A2 => A(2), A3 => A(3), A4 => A(0), ZN 
                           => n28);
   U26 : NAND2_X1 port map( A1 => n25, A2 => n26, ZN => n18);
   U27 : NOR2_X1 port map( A1 => n49, A2 => n50, ZN => n48);
   U28 : XOR2_X1 port map( A => n23, B => A(18), Z => SUM_18_port);
   U29 : XOR2_X1 port map( A => n22, B => A(10), Z => SUM_10_port);
   U30 : OR2_X1 port map( A1 => n70, A2 => n71, ZN => n19);
   U31 : NOR2_X1 port map( A1 => n74, A2 => n75, ZN => n73);
   U32 : XNOR2_X1 port map( A => A(14), B => n67, ZN => SUM_14_port);
   U33 : XNOR2_X1 port map( A => n18, B => A(24), ZN => SUM_24_port);
   U34 : XNOR2_X1 port map( A => n6, B => n38, ZN => SUM_2_port);
   U35 : XNOR2_X1 port map( A => A(17), B => n61, ZN => SUM_17_port);
   U36 : XNOR2_X1 port map( A => A(21), B => n54, ZN => SUM_21_port);
   U37 : NAND2_X1 port map( A1 => A(20), A2 => n55, ZN => n54);
   U38 : XNOR2_X1 port map( A => A(13), B => n69, ZN => SUM_13_port);
   U39 : NAND2_X1 port map( A1 => A(12), A2 => n2, ZN => n69);
   U40 : XNOR2_X1 port map( A => n10, B => n35, ZN => SUM_5_port);
   U41 : XNOR2_X1 port map( A => n20, B => A(26), ZN => SUM_26_port);
   U42 : NAND3_X1 port map( A1 => A(24), A2 => A(25), A3 => n11, ZN => n20);
   U43 : XOR2_X1 port map( A => n44, B => A(29), Z => SUM_29_port);
   U44 : NOR2_X1 port map( A1 => n64, A2 => n65, ZN => n63);
   U45 : XOR2_X1 port map( A => A(27), B => n21, Z => SUM_27_port);
   U46 : AND2_X1 port map( A1 => n27, A2 => A(26), ZN => n21);
   U47 : XNOR2_X1 port map( A => A(6), B => n34, ZN => SUM_6_port);
   U48 : XOR2_X1 port map( A => n16, B => n17, Z => SUM_4_port);
   U49 : XOR2_X1 port map( A => n42, B => A(30), Z => SUM_30_port);
   U50 : XOR2_X1 port map( A => n39, B => A(31), Z => SUM_31_port);
   U51 : XNOR2_X1 port map( A => A(9), B => n29, ZN => SUM_9_port);
   U52 : NAND2_X1 port map( A1 => A(8), A2 => n30, ZN => n29);
   U53 : XNOR2_X1 port map( A => A(3), B => n36, ZN => SUM_3_port);
   U54 : NAND2_X1 port map( A1 => n6, A2 => n37, ZN => n36);
   U55 : INV_X1 port map( A => n38, ZN => n37);
   U56 : AND3_X1 port map( A1 => A(8), A2 => A(9), A3 => n30, ZN => n22);
   U57 : AND3_X1 port map( A1 => A(16), A2 => A(17), A3 => n62, ZN => n23);
   U58 : INV_X1 port map( A => A(28), ZN => n45);
   U59 : NAND2_X1 port map( A1 => A(16), A2 => n62, ZN => n61);
   U60 : NAND2_X1 port map( A1 => n62, A2 => n56, ZN => n53);
   U61 : XNOR2_X1 port map( A => A(22), B => n52, ZN => SUM_22_port);
   U62 : XOR2_X1 port map( A => A(23), B => n24, Z => SUM_23_port);
   U63 : AND2_X1 port map( A1 => n51, A2 => A(22), ZN => n24);
   U64 : AND2_X1 port map( A1 => n48, A2 => n56, ZN => n26);
   U65 : XNOR2_X1 port map( A => A(28), B => n41, ZN => SUM_28_port);
   U66 : NOR2_X1 port map( A1 => n41, A2 => n45, ZN => n44);
   U67 : NOR2_X1 port map( A1 => n41, A2 => n43, ZN => n42);
   U68 : NOR2_X1 port map( A1 => n40, A2 => n41, ZN => n39);
   U69 : NAND2_X1 port map( A1 => n15, A2 => n63, ZN => n60);
   U70 : AND3_X1 port map( A1 => A(24), A2 => A(25), A3 => n11, ZN => n27);
   U71 : NOR2_X1 port map( A1 => n57, A2 => n58, ZN => n56);
   U72 : XNOR2_X1 port map( A => n60, B => A(16), ZN => SUM_16_port);
   U73 : XNOR2_X1 port map( A => A(12), B => n68, ZN => SUM_12_port);
   U74 : INV_X1 port map( A => n60, ZN => n62);
   U75 : XNOR2_X1 port map( A => A(20), B => n53, ZN => SUM_20_port);
   U76 : XNOR2_X1 port map( A => A(8), B => n9, ZN => SUM_8_port);
   U77 : INV_X1 port map( A => n53, ZN => n55);
   U78 : INV_X1 port map( A => n31, ZN => n30);
   U79 : NAND2_X1 port map( A1 => n16, A2 => n17, ZN => n35);
   U80 : NAND2_X1 port map( A1 => n73, A2 => n28, ZN => n31);
   U81 : INV_X1 port map( A => A(0), ZN => SUM_0_port);
   U82 : NAND2_X1 port map( A1 => A(1), A2 => n13, ZN => n38);
   U83 : XNOR2_X1 port map( A => A(7), B => n32, ZN => SUM_7_port);
   U84 : NAND2_X1 port map( A1 => n33, A2 => A(6), ZN => n32);
   U85 : INV_X1 port map( A => n34, ZN => n33);
   U86 : NAND3_X1 port map( A1 => A(4), A2 => n10, A3 => n17, ZN => n34);
   U87 : NAND3_X1 port map( A1 => A(30), A2 => A(29), A3 => A(28), ZN => n40);
   U88 : NAND2_X1 port map( A1 => A(28), A2 => A(29), ZN => n43);
   U89 : NAND2_X1 port map( A1 => A(24), A2 => A(25), ZN => n47);
   U90 : NAND2_X1 port map( A1 => A(27), A2 => A(26), ZN => n46);
   U91 : NAND2_X1 port map( A1 => A(20), A2 => A(21), ZN => n50);
   U92 : NAND2_X1 port map( A1 => A(23), A2 => A(22), ZN => n49);
   U93 : NAND3_X1 port map( A1 => A(20), A2 => A(21), A3 => n55, ZN => n52);
   U94 : NAND2_X1 port map( A1 => A(16), A2 => A(17), ZN => n58);
   U95 : NAND2_X1 port map( A1 => A(19), A2 => A(18), ZN => n57);
   U96 : XOR2_X1 port map( A => A(1), B => n13, Z => SUM_1_port);
   U97 : XNOR2_X1 port map( A => A(19), B => n59, ZN => SUM_19_port);
   U98 : NAND2_X1 port map( A1 => n23, A2 => A(18), ZN => n59);
   U99 : NAND2_X1 port map( A1 => A(12), A2 => A(13), ZN => n65);
   U100 : NAND2_X1 port map( A1 => A(15), A2 => A(14), ZN => n64);
   U101 : INV_X1 port map( A => n67, ZN => n66);
   U102 : NAND3_X1 port map( A1 => A(12), A2 => A(13), A3 => n14, ZN => n67);
   U103 : NAND2_X1 port map( A1 => A(8), A2 => A(9), ZN => n71);
   U104 : NAND2_X1 port map( A1 => A(11), A2 => A(10), ZN => n70);
   U105 : XNOR2_X1 port map( A => A(11), B => n72, ZN => SUM_11_port);
   U106 : NAND2_X1 port map( A1 => n22, A2 => A(10), ZN => n72);
   U107 : NAND2_X1 port map( A1 => A(4), A2 => A(5), ZN => n75);
   U108 : NAND2_X1 port map( A1 => A(7), A2 => A(6), ZN => n74);

end SYN_cla;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity 
   dlx_cu_MICROCODE_MEM_SIZE62_FUNC_SIZE11_OP_CODE_SIZE6_IR_SIZE32_CW_SIZE15_DW01_inc_3 
   is

   port( A : in std_logic_vector (31 downto 0);  SUM : out std_logic_vector (31
         downto 0));

end 
   dlx_cu_MICROCODE_MEM_SIZE62_FUNC_SIZE11_OP_CODE_SIZE6_IR_SIZE32_CW_SIZE15_DW01_inc_3;

architecture SYN_cla of 
   dlx_cu_MICROCODE_MEM_SIZE62_FUNC_SIZE11_OP_CODE_SIZE6_IR_SIZE32_CW_SIZE15_DW01_inc_3 
   is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      , n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, 
      n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45
      , n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, 
      n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74
      , n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, 
      n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, 
      n103, n104, n105, n106 : std_logic;

begin
   
   U2 : CLKBUF_X1 port map( A => A(7), Z => n1);
   U3 : NAND2_X1 port map( A1 => A(7), A2 => A(6), ZN => n2);
   U4 : AND2_X1 port map( A1 => n69, A2 => n37, ZN => n28);
   U5 : AND2_X1 port map( A1 => n69, A2 => n6, ZN => n57);
   U6 : BUF_X1 port map( A => A(1), Z => n8);
   U7 : AND2_X1 port map( A1 => A(12), A2 => n21, ZN => n3);
   U8 : AND2_X1 port map( A1 => A(20), A2 => A(21), ZN => n4);
   U9 : AND2_X1 port map( A1 => A(24), A2 => A(25), ZN => n5);
   U10 : NOR2_X1 port map( A1 => n85, A2 => n86, ZN => n6);
   U11 : XOR2_X1 port map( A => A(22), B => n7, Z => SUM(22));
   U12 : AND2_X1 port map( A1 => n88, A2 => n4, ZN => n7);
   U13 : NOR2_X1 port map( A1 => n65, A2 => n2, ZN => n9);
   U14 : CLKBUF_X1 port map( A => A(0), Z => n10);
   U15 : INV_X1 port map( A => n87, ZN => n11);
   U16 : CLKBUF_X1 port map( A => A(11), Z => n12);
   U17 : INV_X1 port map( A => n74, ZN => n13);
   U18 : CLKBUF_X1 port map( A => n92, Z => n14);
   U19 : CLKBUF_X1 port map( A => A(9), Z => n15);
   U20 : CLKBUF_X1 port map( A => A(10), Z => n16);
   U21 : XNOR2_X1 port map( A => n81, B => n17, ZN => SUM(28));
   U22 : NOR2_X1 port map( A1 => n27, A2 => n59, ZN => n17);
   U23 : INV_X1 port map( A => A(28), ZN => n81);
   U24 : XOR2_X1 port map( A => A(21), B => n18, Z => SUM(21));
   U25 : AND2_X1 port map( A1 => n88, A2 => A(20), ZN => n18);
   U26 : XOR2_X1 port map( A => A(25), B => n19, Z => SUM(25));
   U27 : AND2_X1 port map( A1 => A(24), A2 => n44, ZN => n19);
   U28 : CLKBUF_X1 port map( A => A(15), Z => n20);
   U29 : CLKBUF_X1 port map( A => A(13), Z => n21);
   U30 : AND2_X1 port map( A1 => n53, A2 => n3, ZN => n22);
   U31 : XOR2_X1 port map( A => n1, B => n23, Z => SUM(7));
   U32 : AND2_X1 port map( A1 => n70, A2 => n45, ZN => n23);
   U33 : BUF_X1 port map( A => A(3), Z => n34);
   U34 : XOR2_X1 port map( A => A(26), B => n24, Z => SUM(26));
   U35 : AND2_X1 port map( A1 => n44, A2 => n5, ZN => n24);
   U36 : CLKBUF_X1 port map( A => A(8), Z => n25);
   U37 : BUF_X1 port map( A => A(2), Z => n40);
   U38 : NAND4_X1 port map( A1 => A(15), A2 => A(13), A3 => A(12), A4 => A(14),
                           ZN => n26);
   U39 : INV_X1 port map( A => n28, ZN => n93);
   U40 : NAND2_X1 port map( A1 => n57, A2 => n56, ZN => n27);
   U41 : AND2_X1 port map( A1 => n5, A2 => A(26), ZN => n29);
   U42 : XOR2_X1 port map( A => A(27), B => n30, Z => SUM(27));
   U43 : AND2_X1 port map( A1 => n44, A2 => n29, ZN => n30);
   U44 : NAND4_X1 port map( A1 => A(9), A2 => A(10), A3 => A(11), A4 => A(8), 
                           ZN => n31);
   U45 : NOR2_X1 port map( A1 => n27, A2 => n32, ZN => n78);
   U46 : OR2_X1 port map( A1 => n59, A2 => n79, ZN => n32);
   U47 : CLKBUF_X1 port map( A => n10, Z => n33);
   U48 : AND2_X1 port map( A1 => n35, A2 => n36, ZN => n80);
   U49 : NOR2_X1 port map( A1 => n84, A2 => n59, ZN => n35);
   U50 : AND2_X1 port map( A1 => A(28), A2 => A(29), ZN => n36);
   U51 : AND2_X1 port map( A1 => n102, A2 => n103, ZN => n69);
   U52 : NOR2_X1 port map( A1 => n31, A2 => n26, ZN => n37);
   U53 : OR2_X1 port map( A1 => n81, A2 => n59, ZN => n38);
   U54 : XOR2_X1 port map( A => A(19), B => n39, Z => SUM(19));
   U55 : AND2_X1 port map( A1 => n91, A2 => A(18), ZN => n39);
   U56 : CLKBUF_X1 port map( A => A(5), Z => n41);
   U57 : NAND2_X1 port map( A1 => A(3), A2 => A(2), ZN => n42);
   U58 : NAND2_X1 port map( A1 => n53, A2 => n3, ZN => n97);
   U59 : XOR2_X1 port map( A => A(17), B => n43, Z => SUM(17));
   U60 : AND2_X1 port map( A1 => n28, A2 => A(16), ZN => n43);
   U61 : AND2_X1 port map( A1 => n57, A2 => n56, ZN => n44);
   U62 : CLKBUF_X1 port map( A => A(6), Z => n45);
   U63 : AND2_X1 port map( A1 => n11, A2 => n4, ZN => n46);
   U64 : CLKBUF_X1 port map( A => A(14), Z => n47);
   U65 : CLKBUF_X1 port map( A => A(4), Z => n48);
   U66 : CLKBUF_X1 port map( A => A(12), Z => n49);
   U67 : CLKBUF_X1 port map( A => n67, Z => n50);
   U68 : INV_X1 port map( A => n53, ZN => n99);
   U69 : AND2_X1 port map( A1 => n9, A2 => n68, ZN => n67);
   U70 : CLKBUF_X1 port map( A => n104, Z => n51);
   U71 : CLKBUF_X1 port map( A => n25, Z => n52);
   U72 : AND2_X2 port map( A1 => n67, A2 => n55, ZN => n53);
   U73 : NOR2_X1 port map( A1 => n89, A2 => n90, ZN => n54);
   U74 : AND4_X1 port map( A1 => n12, A2 => A(10), A3 => A(9), A4 => n25, ZN =>
                           n55);
   U75 : AND2_X1 port map( A1 => n54, A2 => n37, ZN => n56);
   U76 : NAND2_X1 port map( A1 => n57, A2 => n56, ZN => n84);
   U77 : NAND2_X1 port map( A1 => n69, A2 => n58, ZN => n87);
   U78 : AND2_X1 port map( A1 => n94, A2 => n54, ZN => n58);
   U79 : OR2_X1 port map( A1 => n82, A2 => n83, ZN => n59);
   U80 : XOR2_X1 port map( A => n20, B => n60, Z => SUM(15));
   U81 : AND2_X1 port map( A1 => n47, A2 => n22, ZN => n60);
   U82 : XOR2_X1 port map( A => n78, B => A(31), Z => SUM(31));
   U83 : XOR2_X1 port map( A => n61, B => A(23), Z => SUM(23));
   U84 : AND2_X1 port map( A1 => n46, A2 => A(22), ZN => n61);
   U85 : XNOR2_X1 port map( A => n47, B => n97, ZN => SUM(14));
   U86 : XNOR2_X1 port map( A => n14, B => A(18), ZN => SUM(18));
   U87 : XNOR2_X1 port map( A => n16, B => n101, ZN => SUM(10));
   U88 : XNOR2_X1 port map( A => n62, B => A(29), ZN => SUM(29));
   U89 : OR2_X1 port map( A1 => n38, A2 => n27, ZN => n62);
   U90 : XOR2_X1 port map( A => n80, B => A(30), Z => SUM(30));
   U91 : XNOR2_X1 port map( A => n49, B => n99, ZN => SUM(12));
   U92 : XOR2_X1 port map( A => n15, B => n63, Z => SUM(9));
   U93 : AND2_X1 port map( A1 => n52, A2 => n50, ZN => n63);
   U94 : XOR2_X1 port map( A => n12, B => n64, Z => SUM(11));
   U95 : AND2_X1 port map( A1 => n100, A2 => n16, ZN => n64);
   U96 : OR2_X1 port map( A1 => n65, A2 => n72, ZN => n71);
   U97 : NAND2_X1 port map( A1 => A(5), A2 => A(4), ZN => n65);
   U98 : XNOR2_X1 port map( A => n41, B => n73, ZN => SUM(5));
   U99 : INV_X1 port map( A => n72, ZN => n74);
   U100 : XOR2_X1 port map( A => n52, B => n50, Z => SUM(8));
   U101 : INV_X1 port map( A => n51, ZN => n76);
   U102 : XNOR2_X1 port map( A => A(24), B => n84, ZN => SUM(24));
   U103 : XNOR2_X1 port map( A => A(16), B => n93, ZN => SUM(16));
   U104 : XNOR2_X1 port map( A => n34, B => n75, ZN => SUM(3));
   U105 : CLKBUF_X1 port map( A => n40, Z => n66);
   U106 : NOR2_X1 port map( A1 => n95, A2 => n96, ZN => n94);
   U107 : NAND4_X1 port map( A1 => A(9), A2 => A(10), A3 => A(11), A4 => A(8), 
                           ZN => n95);
   U108 : NOR2_X1 port map( A1 => n104, A2 => n42, ZN => n68);
   U109 : XNOR2_X1 port map( A => n45, B => n71, ZN => SUM(6));
   U110 : NOR2_X1 port map( A1 => n65, A2 => n106, ZN => n102);
   U111 : NAND2_X1 port map( A1 => n48, A2 => n74, ZN => n73);
   U112 : NOR2_X1 port map( A1 => n77, A2 => n105, ZN => n103);
   U113 : XNOR2_X1 port map( A => n87, B => A(20), ZN => SUM(20));
   U114 : INV_X1 port map( A => n87, ZN => n88);
   U115 : XNOR2_X1 port map( A => n66, B => n51, ZN => SUM(2));
   U116 : NAND2_X1 port map( A1 => n66, A2 => n76, ZN => n75);
   U117 : INV_X1 port map( A => n33, ZN => SUM(0));
   U118 : NAND2_X1 port map( A1 => A(1), A2 => A(0), ZN => n77);
   U119 : NAND4_X1 port map( A1 => n10, A2 => n40, A3 => n8, A4 => n34, ZN => 
                           n72);
   U120 : INV_X1 port map( A => n71, ZN => n70);
   U121 : XNOR2_X1 port map( A => n13, B => n48, ZN => SUM(4));
   U122 : NAND3_X1 port map( A1 => A(30), A2 => A(29), A3 => A(28), ZN => n79);
   U123 : NAND2_X1 port map( A1 => A(24), A2 => A(25), ZN => n83);
   U124 : NAND2_X1 port map( A1 => A(27), A2 => A(26), ZN => n82);
   U125 : NAND2_X1 port map( A1 => A(20), A2 => A(21), ZN => n86);
   U126 : NAND2_X1 port map( A1 => A(23), A2 => A(22), ZN => n85);
   U127 : NAND2_X1 port map( A1 => A(16), A2 => A(17), ZN => n90);
   U128 : NAND2_X1 port map( A1 => A(19), A2 => A(18), ZN => n89);
   U129 : XOR2_X1 port map( A => n8, B => n33, Z => SUM(1));
   U130 : INV_X1 port map( A => n92, ZN => n91);
   U131 : NAND3_X1 port map( A1 => n28, A2 => A(17), A3 => A(16), ZN => n92);
   U132 : NAND4_X1 port map( A1 => A(12), A2 => A(14), A3 => A(13), A4 => A(15)
                           , ZN => n96);
   U133 : XNOR2_X1 port map( A => n21, B => n98, ZN => SUM(13));
   U134 : NAND2_X1 port map( A1 => n53, A2 => n49, ZN => n98);
   U135 : INV_X1 port map( A => n101, ZN => n100);
   U136 : NAND3_X1 port map( A1 => n67, A2 => n15, A3 => n25, ZN => n101);
   U137 : NAND2_X1 port map( A1 => A(3), A2 => A(2), ZN => n105);
   U138 : NAND2_X1 port map( A1 => A(1), A2 => A(0), ZN => n104);
   U139 : NAND2_X1 port map( A1 => A(7), A2 => A(6), ZN => n106);

end SYN_cla;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity windRF_M8_N8_F5_NBIT32_DW01_add_5 is

   port( A, B : in std_logic_vector (6 downto 0);  CI : in std_logic;  SUM : 
         out std_logic_vector (6 downto 0);  CO : out std_logic);

end windRF_M8_N8_F5_NBIT32_DW01_add_5;

architecture SYN_rpl of windRF_M8_N8_F5_NBIT32_DW01_add_5 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal carry_5_port, carry_4_port, carry_3_port, carry_2_port, n4, n5 : 
      std_logic;

begin
   
   U1_4 : FA_X1 port map( A => A(4), B => B(4), CI => carry_4_port, CO => 
                           carry_5_port, S => SUM(4));
   U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => carry_3_port, CO => 
                           carry_4_port, S => SUM(3));
   U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => carry_2_port, CO => 
                           carry_3_port, S => SUM(2));
   U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => n4, CO => carry_2_port, S
                           => SUM(1));
   U1 : XOR2_X1 port map( A => B(0), B => A(0), Z => SUM(0));
   U2 : XNOR2_X1 port map( A => A(6), B => n5, ZN => SUM(6));
   U3 : XOR2_X1 port map( A => A(5), B => carry_5_port, Z => SUM(5));
   U4 : NAND2_X1 port map( A1 => A(5), A2 => carry_5_port, ZN => n5);
   U5 : AND2_X1 port map( A1 => B(0), A2 => A(0), ZN => n4);

end SYN_rpl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity windRF_M8_N8_F5_NBIT32_DW01_add_3 is

   port( A, B : in std_logic_vector (6 downto 0);  CI : in std_logic;  SUM : 
         out std_logic_vector (6 downto 0);  CO : out std_logic);

end windRF_M8_N8_F5_NBIT32_DW01_add_3;

architecture SYN_rpl of windRF_M8_N8_F5_NBIT32_DW01_add_3 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal carry_5_port, carry_4_port, carry_3_port, carry_2_port, n4, n5 : 
      std_logic;

begin
   
   U1_4 : FA_X1 port map( A => A(4), B => B(4), CI => carry_4_port, CO => 
                           carry_5_port, S => SUM(4));
   U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => carry_3_port, CO => 
                           carry_4_port, S => SUM(3));
   U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => carry_2_port, CO => 
                           carry_3_port, S => SUM(2));
   U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => n4, CO => carry_2_port, S
                           => SUM(1));
   U1 : XOR2_X1 port map( A => A(5), B => carry_5_port, Z => SUM(5));
   U2 : XOR2_X1 port map( A => B(0), B => A(0), Z => SUM(0));
   U3 : XNOR2_X1 port map( A => A(6), B => n5, ZN => SUM(6));
   U4 : NAND2_X1 port map( A1 => A(5), A2 => carry_5_port, ZN => n5);
   U5 : AND2_X1 port map( A1 => B(0), A2 => A(0), ZN => n4);

end SYN_rpl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity windRF_M8_N8_F5_NBIT32_DW01_add_1 is

   port( A, B : in std_logic_vector (6 downto 0);  CI : in std_logic;  SUM : 
         out std_logic_vector (6 downto 0);  CO : out std_logic);

end windRF_M8_N8_F5_NBIT32_DW01_add_1;

architecture SYN_rpl of windRF_M8_N8_F5_NBIT32_DW01_add_1 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal carry_5_port, carry_4_port, carry_3_port, carry_2_port, n4, n5 : 
      std_logic;

begin
   
   U1_4 : FA_X1 port map( A => A(4), B => B(4), CI => carry_4_port, CO => 
                           carry_5_port, S => SUM(4));
   U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => carry_3_port, CO => 
                           carry_4_port, S => SUM(3));
   U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => carry_2_port, CO => 
                           carry_3_port, S => SUM(2));
   U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => n4, CO => carry_2_port, S
                           => SUM(1));
   U1 : XOR2_X1 port map( A => A(5), B => carry_5_port, Z => SUM(5));
   U2 : XOR2_X1 port map( A => B(0), B => A(0), Z => SUM(0));
   U3 : XNOR2_X1 port map( A => A(6), B => n5, ZN => SUM(6));
   U4 : NAND2_X1 port map( A1 => A(5), A2 => carry_5_port, ZN => n5);
   U5 : AND2_X1 port map( A1 => B(0), A2 => A(0), ZN => n4);

end SYN_rpl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity SHIFTER_GENERIC_N32_DW_rbsh_0 is

   port( A : in std_logic_vector (31 downto 0);  SH : in std_logic_vector (4 
         downto 0);  SH_TC : in std_logic;  B : out std_logic_vector (31 downto
         0));

end SHIFTER_GENERIC_N32_DW_rbsh_0;

architecture SYN_mx2 of SHIFTER_GENERIC_N32_DW_rbsh_0 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   signal MR_int_1_31_port, MR_int_1_30_port, MR_int_1_29_port, 
      MR_int_1_28_port, MR_int_1_27_port, MR_int_1_26_port, MR_int_1_25_port, 
      MR_int_1_24_port, MR_int_1_23_port, MR_int_1_22_port, MR_int_1_21_port, 
      MR_int_1_20_port, MR_int_1_19_port, MR_int_1_18_port, MR_int_1_17_port, 
      MR_int_1_16_port, MR_int_1_15_port, MR_int_1_14_port, MR_int_1_13_port, 
      MR_int_1_12_port, MR_int_1_11_port, MR_int_1_10_port, MR_int_1_9_port, 
      MR_int_1_8_port, MR_int_1_7_port, MR_int_1_6_port, MR_int_1_5_port, 
      MR_int_1_4_port, MR_int_1_3_port, MR_int_1_2_port, MR_int_1_1_port, 
      MR_int_1_0_port, MR_int_2_31_port, MR_int_2_30_port, MR_int_2_29_port, 
      MR_int_2_28_port, MR_int_2_27_port, MR_int_2_26_port, MR_int_2_25_port, 
      MR_int_2_24_port, MR_int_2_23_port, MR_int_2_22_port, MR_int_2_21_port, 
      MR_int_2_20_port, MR_int_2_19_port, MR_int_2_18_port, MR_int_2_17_port, 
      MR_int_2_16_port, MR_int_2_15_port, MR_int_2_14_port, MR_int_2_13_port, 
      MR_int_2_12_port, MR_int_2_11_port, MR_int_2_10_port, MR_int_2_9_port, 
      MR_int_2_8_port, MR_int_2_7_port, MR_int_2_6_port, MR_int_2_5_port, 
      MR_int_2_4_port, MR_int_2_3_port, MR_int_2_2_port, MR_int_2_1_port, 
      MR_int_2_0_port, MR_int_3_31_port, MR_int_3_30_port, MR_int_3_29_port, 
      MR_int_3_28_port, MR_int_3_27_port, MR_int_3_26_port, MR_int_3_25_port, 
      MR_int_3_24_port, MR_int_3_23_port, MR_int_3_22_port, MR_int_3_21_port, 
      MR_int_3_20_port, MR_int_3_19_port, MR_int_3_18_port, MR_int_3_17_port, 
      MR_int_3_16_port, MR_int_3_15_port, MR_int_3_14_port, MR_int_3_13_port, 
      MR_int_3_12_port, MR_int_3_11_port, MR_int_3_10_port, MR_int_3_9_port, 
      MR_int_3_8_port, MR_int_3_7_port, MR_int_3_6_port, MR_int_3_5_port, 
      MR_int_3_4_port, MR_int_3_3_port, MR_int_3_2_port, MR_int_3_1_port, 
      MR_int_3_0_port, MR_int_4_31_port, MR_int_4_30_port, MR_int_4_29_port, 
      MR_int_4_28_port, MR_int_4_27_port, MR_int_4_26_port, MR_int_4_25_port, 
      MR_int_4_24_port, MR_int_4_23_port, MR_int_4_22_port, MR_int_4_21_port, 
      MR_int_4_20_port, MR_int_4_19_port, MR_int_4_18_port, MR_int_4_17_port, 
      MR_int_4_16_port, MR_int_4_15_port, MR_int_4_14_port, MR_int_4_13_port, 
      MR_int_4_12_port, MR_int_4_11_port, MR_int_4_10_port, MR_int_4_9_port, 
      MR_int_4_8_port, MR_int_4_7_port, MR_int_4_6_port, MR_int_4_5_port, 
      MR_int_4_4_port, MR_int_4_3_port, MR_int_4_2_port, MR_int_4_1_port, 
      MR_int_4_0_port, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, 
      n14, n15 : std_logic;

begin
   
   M1_4_31 : MUX2_X1 port map( A => MR_int_4_31_port, B => MR_int_4_15_port, S 
                           => n15, Z => B(31));
   M1_4_30 : MUX2_X1 port map( A => MR_int_4_30_port, B => MR_int_4_14_port, S 
                           => n15, Z => B(30));
   M1_4_29 : MUX2_X1 port map( A => MR_int_4_29_port, B => MR_int_4_13_port, S 
                           => n15, Z => B(29));
   M1_4_28 : MUX2_X1 port map( A => MR_int_4_28_port, B => MR_int_4_12_port, S 
                           => n15, Z => B(28));
   M1_4_27 : MUX2_X1 port map( A => MR_int_4_27_port, B => MR_int_4_11_port, S 
                           => n15, Z => B(27));
   M1_4_26 : MUX2_X1 port map( A => MR_int_4_26_port, B => MR_int_4_10_port, S 
                           => n15, Z => B(26));
   M1_4_25 : MUX2_X1 port map( A => MR_int_4_25_port, B => MR_int_4_9_port, S 
                           => n15, Z => B(25));
   M1_4_24 : MUX2_X1 port map( A => MR_int_4_24_port, B => MR_int_4_8_port, S 
                           => n15, Z => B(24));
   M1_4_23 : MUX2_X1 port map( A => MR_int_4_23_port, B => MR_int_4_7_port, S 
                           => n14, Z => B(23));
   M1_4_22 : MUX2_X1 port map( A => MR_int_4_22_port, B => MR_int_4_6_port, S 
                           => n14, Z => B(22));
   M1_4_21 : MUX2_X1 port map( A => MR_int_4_21_port, B => MR_int_4_5_port, S 
                           => n14, Z => B(21));
   M1_4_20 : MUX2_X1 port map( A => MR_int_4_20_port, B => MR_int_4_4_port, S 
                           => n14, Z => B(20));
   M1_4_19 : MUX2_X1 port map( A => MR_int_4_19_port, B => MR_int_4_3_port, S 
                           => n14, Z => B(19));
   M1_4_18 : MUX2_X1 port map( A => MR_int_4_18_port, B => MR_int_4_2_port, S 
                           => n14, Z => B(18));
   M1_4_17 : MUX2_X1 port map( A => MR_int_4_17_port, B => MR_int_4_1_port, S 
                           => n14, Z => B(17));
   M1_4_16 : MUX2_X1 port map( A => MR_int_4_16_port, B => MR_int_4_0_port, S 
                           => n14, Z => B(16));
   M1_4_15 : MUX2_X1 port map( A => MR_int_4_15_port, B => MR_int_4_31_port, S 
                           => n14, Z => B(15));
   M1_4_14 : MUX2_X1 port map( A => MR_int_4_14_port, B => MR_int_4_30_port, S 
                           => n14, Z => B(14));
   M1_4_13 : MUX2_X1 port map( A => MR_int_4_13_port, B => MR_int_4_29_port, S 
                           => n14, Z => B(13));
   M1_4_12 : MUX2_X1 port map( A => MR_int_4_12_port, B => MR_int_4_28_port, S 
                           => n14, Z => B(12));
   M1_4_11 : MUX2_X1 port map( A => MR_int_4_11_port, B => MR_int_4_27_port, S 
                           => n13, Z => B(11));
   M1_4_10 : MUX2_X1 port map( A => MR_int_4_10_port, B => MR_int_4_26_port, S 
                           => n13, Z => B(10));
   M1_4_9 : MUX2_X1 port map( A => MR_int_4_9_port, B => MR_int_4_25_port, S =>
                           n13, Z => B(9));
   M1_4_8 : MUX2_X1 port map( A => MR_int_4_8_port, B => MR_int_4_24_port, S =>
                           n13, Z => B(8));
   M1_4_7 : MUX2_X1 port map( A => MR_int_4_7_port, B => MR_int_4_23_port, S =>
                           n13, Z => B(7));
   M1_4_6 : MUX2_X1 port map( A => MR_int_4_6_port, B => MR_int_4_22_port, S =>
                           n13, Z => B(6));
   M1_4_5 : MUX2_X1 port map( A => MR_int_4_5_port, B => MR_int_4_21_port, S =>
                           n13, Z => B(5));
   M1_4_4 : MUX2_X1 port map( A => MR_int_4_4_port, B => MR_int_4_20_port, S =>
                           n13, Z => B(4));
   M1_4_3 : MUX2_X1 port map( A => MR_int_4_3_port, B => MR_int_4_19_port, S =>
                           n13, Z => B(3));
   M1_4_2 : MUX2_X1 port map( A => MR_int_4_2_port, B => MR_int_4_18_port, S =>
                           n13, Z => B(2));
   M1_4_1 : MUX2_X1 port map( A => MR_int_4_1_port, B => MR_int_4_17_port, S =>
                           n13, Z => B(1));
   M1_4_0 : MUX2_X1 port map( A => MR_int_4_0_port, B => MR_int_4_16_port, S =>
                           n13, Z => B(0));
   M1_3_31_0 : MUX2_X1 port map( A => MR_int_3_31_port, B => MR_int_3_7_port, S
                           => n12, Z => MR_int_4_31_port);
   M1_3_30_0 : MUX2_X1 port map( A => MR_int_3_30_port, B => MR_int_3_6_port, S
                           => n12, Z => MR_int_4_30_port);
   M1_3_29_0 : MUX2_X1 port map( A => MR_int_3_29_port, B => MR_int_3_5_port, S
                           => n12, Z => MR_int_4_29_port);
   M1_3_28_0 : MUX2_X1 port map( A => MR_int_3_28_port, B => MR_int_3_4_port, S
                           => n12, Z => MR_int_4_28_port);
   M1_3_27_0 : MUX2_X1 port map( A => MR_int_3_27_port, B => MR_int_3_3_port, S
                           => n12, Z => MR_int_4_27_port);
   M1_3_26_0 : MUX2_X1 port map( A => MR_int_3_26_port, B => MR_int_3_2_port, S
                           => n12, Z => MR_int_4_26_port);
   M1_3_25_0 : MUX2_X1 port map( A => MR_int_3_25_port, B => MR_int_3_1_port, S
                           => n12, Z => MR_int_4_25_port);
   M1_3_24_0 : MUX2_X1 port map( A => MR_int_3_24_port, B => MR_int_3_0_port, S
                           => n12, Z => MR_int_4_24_port);
   M1_3_23_0 : MUX2_X1 port map( A => MR_int_3_23_port, B => MR_int_3_31_port, 
                           S => n11, Z => MR_int_4_23_port);
   M1_3_22_0 : MUX2_X1 port map( A => MR_int_3_22_port, B => MR_int_3_30_port, 
                           S => n11, Z => MR_int_4_22_port);
   M1_3_21_0 : MUX2_X1 port map( A => MR_int_3_21_port, B => MR_int_3_29_port, 
                           S => n11, Z => MR_int_4_21_port);
   M1_3_20_0 : MUX2_X1 port map( A => MR_int_3_20_port, B => MR_int_3_28_port, 
                           S => n11, Z => MR_int_4_20_port);
   M1_3_19_0 : MUX2_X1 port map( A => MR_int_3_19_port, B => MR_int_3_27_port, 
                           S => n11, Z => MR_int_4_19_port);
   M1_3_18_0 : MUX2_X1 port map( A => MR_int_3_18_port, B => MR_int_3_26_port, 
                           S => n11, Z => MR_int_4_18_port);
   M1_3_17_0 : MUX2_X1 port map( A => MR_int_3_17_port, B => MR_int_3_25_port, 
                           S => n11, Z => MR_int_4_17_port);
   M1_3_16_0 : MUX2_X1 port map( A => MR_int_3_16_port, B => MR_int_3_24_port, 
                           S => n11, Z => MR_int_4_16_port);
   M1_3_15_0 : MUX2_X1 port map( A => MR_int_3_15_port, B => MR_int_3_23_port, 
                           S => n11, Z => MR_int_4_15_port);
   M1_3_14_0 : MUX2_X1 port map( A => MR_int_3_14_port, B => MR_int_3_22_port, 
                           S => n11, Z => MR_int_4_14_port);
   M1_3_13_0 : MUX2_X1 port map( A => MR_int_3_13_port, B => MR_int_3_21_port, 
                           S => n11, Z => MR_int_4_13_port);
   M1_3_12_0 : MUX2_X1 port map( A => MR_int_3_12_port, B => MR_int_3_20_port, 
                           S => n11, Z => MR_int_4_12_port);
   M1_3_11_0 : MUX2_X1 port map( A => MR_int_3_11_port, B => MR_int_3_19_port, 
                           S => n10, Z => MR_int_4_11_port);
   M1_3_10_0 : MUX2_X1 port map( A => MR_int_3_10_port, B => MR_int_3_18_port, 
                           S => n10, Z => MR_int_4_10_port);
   M1_3_9_0 : MUX2_X1 port map( A => MR_int_3_9_port, B => MR_int_3_17_port, S 
                           => n10, Z => MR_int_4_9_port);
   M1_3_8_0 : MUX2_X1 port map( A => MR_int_3_8_port, B => MR_int_3_16_port, S 
                           => n10, Z => MR_int_4_8_port);
   M1_3_7 : MUX2_X1 port map( A => MR_int_3_7_port, B => MR_int_3_15_port, S =>
                           n10, Z => MR_int_4_7_port);
   M1_3_6 : MUX2_X1 port map( A => MR_int_3_6_port, B => MR_int_3_14_port, S =>
                           n10, Z => MR_int_4_6_port);
   M1_3_5 : MUX2_X1 port map( A => MR_int_3_5_port, B => MR_int_3_13_port, S =>
                           n10, Z => MR_int_4_5_port);
   M1_3_4 : MUX2_X1 port map( A => MR_int_3_4_port, B => MR_int_3_12_port, S =>
                           n10, Z => MR_int_4_4_port);
   M1_3_3 : MUX2_X1 port map( A => MR_int_3_3_port, B => MR_int_3_11_port, S =>
                           n10, Z => MR_int_4_3_port);
   M1_3_2 : MUX2_X1 port map( A => MR_int_3_2_port, B => MR_int_3_10_port, S =>
                           n10, Z => MR_int_4_2_port);
   M1_3_1 : MUX2_X1 port map( A => MR_int_3_1_port, B => MR_int_3_9_port, S => 
                           n10, Z => MR_int_4_1_port);
   M1_3_0 : MUX2_X1 port map( A => MR_int_3_0_port, B => MR_int_3_8_port, S => 
                           n10, Z => MR_int_4_0_port);
   M1_2_31_0 : MUX2_X1 port map( A => MR_int_2_31_port, B => MR_int_2_3_port, S
                           => n9, Z => MR_int_3_31_port);
   M1_2_30_0 : MUX2_X1 port map( A => MR_int_2_30_port, B => MR_int_2_2_port, S
                           => n9, Z => MR_int_3_30_port);
   M1_2_29_0 : MUX2_X1 port map( A => MR_int_2_29_port, B => MR_int_2_1_port, S
                           => n9, Z => MR_int_3_29_port);
   M1_2_28_0 : MUX2_X1 port map( A => MR_int_2_28_port, B => MR_int_2_0_port, S
                           => n9, Z => MR_int_3_28_port);
   M1_2_27_0 : MUX2_X1 port map( A => MR_int_2_27_port, B => MR_int_2_31_port, 
                           S => n9, Z => MR_int_3_27_port);
   M1_2_26_0 : MUX2_X1 port map( A => MR_int_2_26_port, B => MR_int_2_30_port, 
                           S => n9, Z => MR_int_3_26_port);
   M1_2_25_0 : MUX2_X1 port map( A => MR_int_2_25_port, B => MR_int_2_29_port, 
                           S => n9, Z => MR_int_3_25_port);
   M1_2_24_0 : MUX2_X1 port map( A => MR_int_2_24_port, B => MR_int_2_28_port, 
                           S => n9, Z => MR_int_3_24_port);
   M1_2_23_0 : MUX2_X1 port map( A => MR_int_2_23_port, B => MR_int_2_27_port, 
                           S => n8, Z => MR_int_3_23_port);
   M1_2_22_0 : MUX2_X1 port map( A => MR_int_2_22_port, B => MR_int_2_26_port, 
                           S => n8, Z => MR_int_3_22_port);
   M1_2_21_0 : MUX2_X1 port map( A => MR_int_2_21_port, B => MR_int_2_25_port, 
                           S => n8, Z => MR_int_3_21_port);
   M1_2_20_0 : MUX2_X1 port map( A => MR_int_2_20_port, B => MR_int_2_24_port, 
                           S => n8, Z => MR_int_3_20_port);
   M1_2_19_0 : MUX2_X1 port map( A => MR_int_2_19_port, B => MR_int_2_23_port, 
                           S => n8, Z => MR_int_3_19_port);
   M1_2_18_0 : MUX2_X1 port map( A => MR_int_2_18_port, B => MR_int_2_22_port, 
                           S => n8, Z => MR_int_3_18_port);
   M1_2_17_0 : MUX2_X1 port map( A => MR_int_2_17_port, B => MR_int_2_21_port, 
                           S => n8, Z => MR_int_3_17_port);
   M1_2_16_0 : MUX2_X1 port map( A => MR_int_2_16_port, B => MR_int_2_20_port, 
                           S => n8, Z => MR_int_3_16_port);
   M1_2_15_0 : MUX2_X1 port map( A => MR_int_2_15_port, B => MR_int_2_19_port, 
                           S => n8, Z => MR_int_3_15_port);
   M1_2_14_0 : MUX2_X1 port map( A => MR_int_2_14_port, B => MR_int_2_18_port, 
                           S => n8, Z => MR_int_3_14_port);
   M1_2_13_0 : MUX2_X1 port map( A => MR_int_2_13_port, B => MR_int_2_17_port, 
                           S => n8, Z => MR_int_3_13_port);
   M1_2_12_0 : MUX2_X1 port map( A => MR_int_2_12_port, B => MR_int_2_16_port, 
                           S => n8, Z => MR_int_3_12_port);
   M1_2_11_0 : MUX2_X1 port map( A => MR_int_2_11_port, B => MR_int_2_15_port, 
                           S => n7, Z => MR_int_3_11_port);
   M1_2_10_0 : MUX2_X1 port map( A => MR_int_2_10_port, B => MR_int_2_14_port, 
                           S => n7, Z => MR_int_3_10_port);
   M1_2_9_0 : MUX2_X1 port map( A => MR_int_2_9_port, B => MR_int_2_13_port, S 
                           => n7, Z => MR_int_3_9_port);
   M1_2_8_0 : MUX2_X1 port map( A => MR_int_2_8_port, B => MR_int_2_12_port, S 
                           => n7, Z => MR_int_3_8_port);
   M1_2_7_0 : MUX2_X1 port map( A => MR_int_2_7_port, B => MR_int_2_11_port, S 
                           => n7, Z => MR_int_3_7_port);
   M1_2_6_0 : MUX2_X1 port map( A => MR_int_2_6_port, B => MR_int_2_10_port, S 
                           => n7, Z => MR_int_3_6_port);
   M1_2_5_0 : MUX2_X1 port map( A => MR_int_2_5_port, B => MR_int_2_9_port, S 
                           => n7, Z => MR_int_3_5_port);
   M1_2_4_0 : MUX2_X1 port map( A => MR_int_2_4_port, B => MR_int_2_8_port, S 
                           => n7, Z => MR_int_3_4_port);
   M1_2_3 : MUX2_X1 port map( A => MR_int_2_3_port, B => MR_int_2_7_port, S => 
                           n7, Z => MR_int_3_3_port);
   M1_2_2 : MUX2_X1 port map( A => MR_int_2_2_port, B => MR_int_2_6_port, S => 
                           n7, Z => MR_int_3_2_port);
   M1_2_1 : MUX2_X1 port map( A => MR_int_2_1_port, B => MR_int_2_5_port, S => 
                           n7, Z => MR_int_3_1_port);
   M1_2_0 : MUX2_X1 port map( A => MR_int_2_0_port, B => MR_int_2_4_port, S => 
                           n7, Z => MR_int_3_0_port);
   M1_1_31_0 : MUX2_X1 port map( A => MR_int_1_31_port, B => MR_int_1_1_port, S
                           => n6, Z => MR_int_2_31_port);
   M1_1_30_0 : MUX2_X1 port map( A => MR_int_1_30_port, B => MR_int_1_0_port, S
                           => n6, Z => MR_int_2_30_port);
   M1_1_29_0 : MUX2_X1 port map( A => MR_int_1_29_port, B => MR_int_1_31_port, 
                           S => n6, Z => MR_int_2_29_port);
   M1_1_28_0 : MUX2_X1 port map( A => MR_int_1_28_port, B => MR_int_1_30_port, 
                           S => n6, Z => MR_int_2_28_port);
   M1_1_27_0 : MUX2_X1 port map( A => MR_int_1_27_port, B => MR_int_1_29_port, 
                           S => n6, Z => MR_int_2_27_port);
   M1_1_26_0 : MUX2_X1 port map( A => MR_int_1_26_port, B => MR_int_1_28_port, 
                           S => n6, Z => MR_int_2_26_port);
   M1_1_25_0 : MUX2_X1 port map( A => MR_int_1_25_port, B => MR_int_1_27_port, 
                           S => n6, Z => MR_int_2_25_port);
   M1_1_24_0 : MUX2_X1 port map( A => MR_int_1_24_port, B => MR_int_1_26_port, 
                           S => n6, Z => MR_int_2_24_port);
   M1_1_23_0 : MUX2_X1 port map( A => MR_int_1_23_port, B => MR_int_1_25_port, 
                           S => n5, Z => MR_int_2_23_port);
   M1_1_22_0 : MUX2_X1 port map( A => MR_int_1_22_port, B => MR_int_1_24_port, 
                           S => n5, Z => MR_int_2_22_port);
   M1_1_21_0 : MUX2_X1 port map( A => MR_int_1_21_port, B => MR_int_1_23_port, 
                           S => n5, Z => MR_int_2_21_port);
   M1_1_20_0 : MUX2_X1 port map( A => MR_int_1_20_port, B => MR_int_1_22_port, 
                           S => n5, Z => MR_int_2_20_port);
   M1_1_19_0 : MUX2_X1 port map( A => MR_int_1_19_port, B => MR_int_1_21_port, 
                           S => n5, Z => MR_int_2_19_port);
   M1_1_18_0 : MUX2_X1 port map( A => MR_int_1_18_port, B => MR_int_1_20_port, 
                           S => n5, Z => MR_int_2_18_port);
   M1_1_17_0 : MUX2_X1 port map( A => MR_int_1_17_port, B => MR_int_1_19_port, 
                           S => n5, Z => MR_int_2_17_port);
   M1_1_16_0 : MUX2_X1 port map( A => MR_int_1_16_port, B => MR_int_1_18_port, 
                           S => n5, Z => MR_int_2_16_port);
   M1_1_15_0 : MUX2_X1 port map( A => MR_int_1_15_port, B => MR_int_1_17_port, 
                           S => n5, Z => MR_int_2_15_port);
   M1_1_14_0 : MUX2_X1 port map( A => MR_int_1_14_port, B => MR_int_1_16_port, 
                           S => n5, Z => MR_int_2_14_port);
   M1_1_13_0 : MUX2_X1 port map( A => MR_int_1_13_port, B => MR_int_1_15_port, 
                           S => n5, Z => MR_int_2_13_port);
   M1_1_12_0 : MUX2_X1 port map( A => MR_int_1_12_port, B => MR_int_1_14_port, 
                           S => n5, Z => MR_int_2_12_port);
   M1_1_11_0 : MUX2_X1 port map( A => MR_int_1_11_port, B => MR_int_1_13_port, 
                           S => n4, Z => MR_int_2_11_port);
   M1_1_10_0 : MUX2_X1 port map( A => MR_int_1_10_port, B => MR_int_1_12_port, 
                           S => n4, Z => MR_int_2_10_port);
   M1_1_9_0 : MUX2_X1 port map( A => MR_int_1_9_port, B => MR_int_1_11_port, S 
                           => n4, Z => MR_int_2_9_port);
   M1_1_8_0 : MUX2_X1 port map( A => MR_int_1_8_port, B => MR_int_1_10_port, S 
                           => n4, Z => MR_int_2_8_port);
   M1_1_7_0 : MUX2_X1 port map( A => MR_int_1_7_port, B => MR_int_1_9_port, S 
                           => n4, Z => MR_int_2_7_port);
   M1_1_6_0 : MUX2_X1 port map( A => MR_int_1_6_port, B => MR_int_1_8_port, S 
                           => n4, Z => MR_int_2_6_port);
   M1_1_5_0 : MUX2_X1 port map( A => MR_int_1_5_port, B => MR_int_1_7_port, S 
                           => n4, Z => MR_int_2_5_port);
   M1_1_4_0 : MUX2_X1 port map( A => MR_int_1_4_port, B => MR_int_1_6_port, S 
                           => n4, Z => MR_int_2_4_port);
   M1_1_3_0 : MUX2_X1 port map( A => MR_int_1_3_port, B => MR_int_1_5_port, S 
                           => n4, Z => MR_int_2_3_port);
   M1_1_2_0 : MUX2_X1 port map( A => MR_int_1_2_port, B => MR_int_1_4_port, S 
                           => n4, Z => MR_int_2_2_port);
   M1_1_1 : MUX2_X1 port map( A => MR_int_1_1_port, B => MR_int_1_3_port, S => 
                           n4, Z => MR_int_2_1_port);
   M1_1_0 : MUX2_X1 port map( A => MR_int_1_0_port, B => MR_int_1_2_port, S => 
                           n4, Z => MR_int_2_0_port);
   M1_0_31_0 : MUX2_X1 port map( A => A(31), B => A(0), S => n3, Z => 
                           MR_int_1_31_port);
   M1_0_30_0 : MUX2_X1 port map( A => A(30), B => A(31), S => n3, Z => 
                           MR_int_1_30_port);
   M1_0_29_0 : MUX2_X1 port map( A => A(29), B => A(30), S => n3, Z => 
                           MR_int_1_29_port);
   M1_0_28_0 : MUX2_X1 port map( A => A(28), B => A(29), S => n3, Z => 
                           MR_int_1_28_port);
   M1_0_27_0 : MUX2_X1 port map( A => A(27), B => A(28), S => n3, Z => 
                           MR_int_1_27_port);
   M1_0_26_0 : MUX2_X1 port map( A => A(26), B => A(27), S => n3, Z => 
                           MR_int_1_26_port);
   M1_0_25_0 : MUX2_X1 port map( A => A(25), B => A(26), S => n3, Z => 
                           MR_int_1_25_port);
   M1_0_24_0 : MUX2_X1 port map( A => A(24), B => A(25), S => n3, Z => 
                           MR_int_1_24_port);
   M1_0_23_0 : MUX2_X1 port map( A => A(23), B => A(24), S => n2, Z => 
                           MR_int_1_23_port);
   M1_0_22_0 : MUX2_X1 port map( A => A(22), B => A(23), S => n2, Z => 
                           MR_int_1_22_port);
   M1_0_21_0 : MUX2_X1 port map( A => A(21), B => A(22), S => n2, Z => 
                           MR_int_1_21_port);
   M1_0_20_0 : MUX2_X1 port map( A => A(20), B => A(21), S => n2, Z => 
                           MR_int_1_20_port);
   M1_0_19_0 : MUX2_X1 port map( A => A(19), B => A(20), S => n2, Z => 
                           MR_int_1_19_port);
   M1_0_18_0 : MUX2_X1 port map( A => A(18), B => A(19), S => n2, Z => 
                           MR_int_1_18_port);
   M1_0_17_0 : MUX2_X1 port map( A => A(17), B => A(18), S => n2, Z => 
                           MR_int_1_17_port);
   M1_0_16_0 : MUX2_X1 port map( A => A(16), B => A(17), S => n2, Z => 
                           MR_int_1_16_port);
   M1_0_15_0 : MUX2_X1 port map( A => A(15), B => A(16), S => n2, Z => 
                           MR_int_1_15_port);
   M1_0_14_0 : MUX2_X1 port map( A => A(14), B => A(15), S => n2, Z => 
                           MR_int_1_14_port);
   M1_0_13_0 : MUX2_X1 port map( A => A(13), B => A(14), S => n2, Z => 
                           MR_int_1_13_port);
   M1_0_12_0 : MUX2_X1 port map( A => A(12), B => A(13), S => n2, Z => 
                           MR_int_1_12_port);
   M1_0_11_0 : MUX2_X1 port map( A => A(11), B => A(12), S => n1, Z => 
                           MR_int_1_11_port);
   M1_0_10_0 : MUX2_X1 port map( A => A(10), B => A(11), S => n1, Z => 
                           MR_int_1_10_port);
   M1_0_9_0 : MUX2_X1 port map( A => A(9), B => A(10), S => n1, Z => 
                           MR_int_1_9_port);
   M1_0_8_0 : MUX2_X1 port map( A => A(8), B => A(9), S => n1, Z => 
                           MR_int_1_8_port);
   M1_0_7_0 : MUX2_X1 port map( A => A(7), B => A(8), S => n1, Z => 
                           MR_int_1_7_port);
   M1_0_6_0 : MUX2_X1 port map( A => A(6), B => A(7), S => n1, Z => 
                           MR_int_1_6_port);
   M1_0_5_0 : MUX2_X1 port map( A => A(5), B => A(6), S => n1, Z => 
                           MR_int_1_5_port);
   M1_0_4_0 : MUX2_X1 port map( A => A(4), B => A(5), S => n1, Z => 
                           MR_int_1_4_port);
   M1_0_3_0 : MUX2_X1 port map( A => A(3), B => A(4), S => n1, Z => 
                           MR_int_1_3_port);
   M1_0_2_0 : MUX2_X1 port map( A => A(2), B => A(3), S => n1, Z => 
                           MR_int_1_2_port);
   M1_0_1_0 : MUX2_X1 port map( A => A(1), B => A(2), S => n1, Z => 
                           MR_int_1_1_port);
   M1_0_0 : MUX2_X1 port map( A => A(0), B => A(1), S => n1, Z => 
                           MR_int_1_0_port);
   U2 : BUF_X1 port map( A => SH(4), Z => n14);
   U3 : BUF_X1 port map( A => SH(4), Z => n13);
   U4 : BUF_X1 port map( A => SH(4), Z => n15);
   U5 : BUF_X1 port map( A => SH(1), Z => n5);
   U6 : BUF_X1 port map( A => SH(1), Z => n4);
   U7 : BUF_X1 port map( A => SH(2), Z => n8);
   U8 : BUF_X1 port map( A => SH(2), Z => n7);
   U9 : BUF_X1 port map( A => SH(0), Z => n2);
   U10 : BUF_X1 port map( A => SH(0), Z => n1);
   U11 : BUF_X1 port map( A => SH(3), Z => n11);
   U12 : BUF_X1 port map( A => SH(3), Z => n10);
   U13 : BUF_X1 port map( A => SH(1), Z => n6);
   U14 : BUF_X1 port map( A => SH(2), Z => n9);
   U15 : BUF_X1 port map( A => SH(0), Z => n3);
   U16 : BUF_X1 port map( A => SH(3), Z => n12);

end SYN_mx2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity SHIFTER_GENERIC_N32_DW_lbsh_0 is

   port( A : in std_logic_vector (31 downto 0);  SH : in std_logic_vector (4 
         downto 0);  SH_TC : in std_logic;  B : out std_logic_vector (31 downto
         0));

end SHIFTER_GENERIC_N32_DW_lbsh_0;

architecture SYN_mx2 of SHIFTER_GENERIC_N32_DW_lbsh_0 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   signal ML_int_1_31_port, ML_int_1_30_port, ML_int_1_29_port, 
      ML_int_1_28_port, ML_int_1_27_port, ML_int_1_26_port, ML_int_1_25_port, 
      ML_int_1_24_port, ML_int_1_23_port, ML_int_1_22_port, ML_int_1_21_port, 
      ML_int_1_20_port, ML_int_1_19_port, ML_int_1_18_port, ML_int_1_17_port, 
      ML_int_1_16_port, ML_int_1_15_port, ML_int_1_14_port, ML_int_1_13_port, 
      ML_int_1_12_port, ML_int_1_11_port, ML_int_1_10_port, ML_int_1_9_port, 
      ML_int_1_8_port, ML_int_1_7_port, ML_int_1_6_port, ML_int_1_5_port, 
      ML_int_1_4_port, ML_int_1_3_port, ML_int_1_2_port, ML_int_1_1_port, 
      ML_int_1_0_port, ML_int_2_31_port, ML_int_2_30_port, ML_int_2_29_port, 
      ML_int_2_28_port, ML_int_2_27_port, ML_int_2_26_port, ML_int_2_25_port, 
      ML_int_2_24_port, ML_int_2_23_port, ML_int_2_22_port, ML_int_2_21_port, 
      ML_int_2_20_port, ML_int_2_19_port, ML_int_2_18_port, ML_int_2_17_port, 
      ML_int_2_16_port, ML_int_2_15_port, ML_int_2_14_port, ML_int_2_13_port, 
      ML_int_2_12_port, ML_int_2_11_port, ML_int_2_10_port, ML_int_2_9_port, 
      ML_int_2_8_port, ML_int_2_7_port, ML_int_2_6_port, ML_int_2_5_port, 
      ML_int_2_4_port, ML_int_2_3_port, ML_int_2_2_port, ML_int_2_1_port, 
      ML_int_2_0_port, ML_int_3_31_port, ML_int_3_30_port, ML_int_3_29_port, 
      ML_int_3_28_port, ML_int_3_27_port, ML_int_3_26_port, ML_int_3_25_port, 
      ML_int_3_24_port, ML_int_3_23_port, ML_int_3_22_port, ML_int_3_21_port, 
      ML_int_3_20_port, ML_int_3_19_port, ML_int_3_18_port, ML_int_3_17_port, 
      ML_int_3_16_port, ML_int_3_15_port, ML_int_3_14_port, ML_int_3_13_port, 
      ML_int_3_12_port, ML_int_3_11_port, ML_int_3_10_port, ML_int_3_9_port, 
      ML_int_3_8_port, ML_int_3_7_port, ML_int_3_6_port, ML_int_3_5_port, 
      ML_int_3_4_port, ML_int_3_3_port, ML_int_3_2_port, ML_int_3_1_port, 
      ML_int_3_0_port, ML_int_4_31_port, ML_int_4_30_port, ML_int_4_29_port, 
      ML_int_4_28_port, ML_int_4_27_port, ML_int_4_26_port, ML_int_4_25_port, 
      ML_int_4_24_port, ML_int_4_23_port, ML_int_4_22_port, ML_int_4_21_port, 
      ML_int_4_20_port, ML_int_4_19_port, ML_int_4_18_port, ML_int_4_17_port, 
      ML_int_4_16_port, ML_int_4_15_port, ML_int_4_14_port, ML_int_4_13_port, 
      ML_int_4_12_port, ML_int_4_11_port, ML_int_4_10_port, ML_int_4_9_port, 
      ML_int_4_8_port, ML_int_4_7_port, ML_int_4_6_port, ML_int_4_5_port, 
      ML_int_4_4_port, ML_int_4_3_port, ML_int_4_2_port, ML_int_4_1_port, 
      ML_int_4_0_port, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, 
      n14, n15 : std_logic;

begin
   
   M1_4_31 : MUX2_X1 port map( A => ML_int_4_31_port, B => ML_int_4_15_port, S 
                           => n15, Z => B(31));
   M1_4_30 : MUX2_X1 port map( A => ML_int_4_30_port, B => ML_int_4_14_port, S 
                           => n15, Z => B(30));
   M1_4_29 : MUX2_X1 port map( A => ML_int_4_29_port, B => ML_int_4_13_port, S 
                           => n15, Z => B(29));
   M1_4_28 : MUX2_X1 port map( A => ML_int_4_28_port, B => ML_int_4_12_port, S 
                           => n15, Z => B(28));
   M1_4_27 : MUX2_X1 port map( A => ML_int_4_27_port, B => ML_int_4_11_port, S 
                           => n15, Z => B(27));
   M1_4_26 : MUX2_X1 port map( A => ML_int_4_26_port, B => ML_int_4_10_port, S 
                           => n15, Z => B(26));
   M1_4_25 : MUX2_X1 port map( A => ML_int_4_25_port, B => ML_int_4_9_port, S 
                           => n15, Z => B(25));
   M1_4_24 : MUX2_X1 port map( A => ML_int_4_24_port, B => ML_int_4_8_port, S 
                           => n15, Z => B(24));
   M1_4_23 : MUX2_X1 port map( A => ML_int_4_23_port, B => ML_int_4_7_port, S 
                           => n14, Z => B(23));
   M1_4_22 : MUX2_X1 port map( A => ML_int_4_22_port, B => ML_int_4_6_port, S 
                           => n14, Z => B(22));
   M1_4_21 : MUX2_X1 port map( A => ML_int_4_21_port, B => ML_int_4_5_port, S 
                           => n14, Z => B(21));
   M1_4_20 : MUX2_X1 port map( A => ML_int_4_20_port, B => ML_int_4_4_port, S 
                           => n14, Z => B(20));
   M1_4_19 : MUX2_X1 port map( A => ML_int_4_19_port, B => ML_int_4_3_port, S 
                           => n14, Z => B(19));
   M1_4_18 : MUX2_X1 port map( A => ML_int_4_18_port, B => ML_int_4_2_port, S 
                           => n14, Z => B(18));
   M1_4_17 : MUX2_X1 port map( A => ML_int_4_17_port, B => ML_int_4_1_port, S 
                           => n14, Z => B(17));
   M1_4_16 : MUX2_X1 port map( A => ML_int_4_16_port, B => ML_int_4_0_port, S 
                           => n14, Z => B(16));
   M0_4_15 : MUX2_X1 port map( A => ML_int_4_15_port, B => ML_int_4_31_port, S 
                           => n14, Z => B(15));
   M0_4_14 : MUX2_X1 port map( A => ML_int_4_14_port, B => ML_int_4_30_port, S 
                           => n14, Z => B(14));
   M0_4_13 : MUX2_X1 port map( A => ML_int_4_13_port, B => ML_int_4_29_port, S 
                           => n14, Z => B(13));
   M0_4_12 : MUX2_X1 port map( A => ML_int_4_12_port, B => ML_int_4_28_port, S 
                           => n14, Z => B(12));
   M0_4_11 : MUX2_X1 port map( A => ML_int_4_11_port, B => ML_int_4_27_port, S 
                           => n13, Z => B(11));
   M0_4_10 : MUX2_X1 port map( A => ML_int_4_10_port, B => ML_int_4_26_port, S 
                           => n13, Z => B(10));
   M0_4_9 : MUX2_X1 port map( A => ML_int_4_9_port, B => ML_int_4_25_port, S =>
                           n13, Z => B(9));
   M0_4_8 : MUX2_X1 port map( A => ML_int_4_8_port, B => ML_int_4_24_port, S =>
                           n13, Z => B(8));
   M0_4_7 : MUX2_X1 port map( A => ML_int_4_7_port, B => ML_int_4_23_port, S =>
                           n13, Z => B(7));
   M0_4_6 : MUX2_X1 port map( A => ML_int_4_6_port, B => ML_int_4_22_port, S =>
                           n13, Z => B(6));
   M0_4_5 : MUX2_X1 port map( A => ML_int_4_5_port, B => ML_int_4_21_port, S =>
                           n13, Z => B(5));
   M0_4_4 : MUX2_X1 port map( A => ML_int_4_4_port, B => ML_int_4_20_port, S =>
                           n13, Z => B(4));
   M0_4_3 : MUX2_X1 port map( A => ML_int_4_3_port, B => ML_int_4_19_port, S =>
                           n13, Z => B(3));
   M0_4_2 : MUX2_X1 port map( A => ML_int_4_2_port, B => ML_int_4_18_port, S =>
                           n13, Z => B(2));
   M0_4_1 : MUX2_X1 port map( A => ML_int_4_1_port, B => ML_int_4_17_port, S =>
                           n13, Z => B(1));
   M0_4_0 : MUX2_X1 port map( A => ML_int_4_0_port, B => ML_int_4_16_port, S =>
                           n13, Z => B(0));
   M1_3_31 : MUX2_X1 port map( A => ML_int_3_31_port, B => ML_int_3_23_port, S 
                           => n12, Z => ML_int_4_31_port);
   M1_3_30 : MUX2_X1 port map( A => ML_int_3_30_port, B => ML_int_3_22_port, S 
                           => n12, Z => ML_int_4_30_port);
   M1_3_29 : MUX2_X1 port map( A => ML_int_3_29_port, B => ML_int_3_21_port, S 
                           => n12, Z => ML_int_4_29_port);
   M1_3_28 : MUX2_X1 port map( A => ML_int_3_28_port, B => ML_int_3_20_port, S 
                           => n12, Z => ML_int_4_28_port);
   M1_3_27 : MUX2_X1 port map( A => ML_int_3_27_port, B => ML_int_3_19_port, S 
                           => n12, Z => ML_int_4_27_port);
   M1_3_26 : MUX2_X1 port map( A => ML_int_3_26_port, B => ML_int_3_18_port, S 
                           => n12, Z => ML_int_4_26_port);
   M1_3_25 : MUX2_X1 port map( A => ML_int_3_25_port, B => ML_int_3_17_port, S 
                           => n12, Z => ML_int_4_25_port);
   M1_3_24 : MUX2_X1 port map( A => ML_int_3_24_port, B => ML_int_3_16_port, S 
                           => n12, Z => ML_int_4_24_port);
   M1_3_23 : MUX2_X1 port map( A => ML_int_3_23_port, B => ML_int_3_15_port, S 
                           => n11, Z => ML_int_4_23_port);
   M1_3_22 : MUX2_X1 port map( A => ML_int_3_22_port, B => ML_int_3_14_port, S 
                           => n11, Z => ML_int_4_22_port);
   M1_3_21 : MUX2_X1 port map( A => ML_int_3_21_port, B => ML_int_3_13_port, S 
                           => n11, Z => ML_int_4_21_port);
   M1_3_20 : MUX2_X1 port map( A => ML_int_3_20_port, B => ML_int_3_12_port, S 
                           => n11, Z => ML_int_4_20_port);
   M1_3_19 : MUX2_X1 port map( A => ML_int_3_19_port, B => ML_int_3_11_port, S 
                           => n11, Z => ML_int_4_19_port);
   M1_3_18 : MUX2_X1 port map( A => ML_int_3_18_port, B => ML_int_3_10_port, S 
                           => n11, Z => ML_int_4_18_port);
   M1_3_17 : MUX2_X1 port map( A => ML_int_3_17_port, B => ML_int_3_9_port, S 
                           => n11, Z => ML_int_4_17_port);
   M1_3_16 : MUX2_X1 port map( A => ML_int_3_16_port, B => ML_int_3_8_port, S 
                           => n11, Z => ML_int_4_16_port);
   M1_3_15 : MUX2_X1 port map( A => ML_int_3_15_port, B => ML_int_3_7_port, S 
                           => n11, Z => ML_int_4_15_port);
   M1_3_14 : MUX2_X1 port map( A => ML_int_3_14_port, B => ML_int_3_6_port, S 
                           => n11, Z => ML_int_4_14_port);
   M1_3_13 : MUX2_X1 port map( A => ML_int_3_13_port, B => ML_int_3_5_port, S 
                           => n11, Z => ML_int_4_13_port);
   M1_3_12 : MUX2_X1 port map( A => ML_int_3_12_port, B => ML_int_3_4_port, S 
                           => n11, Z => ML_int_4_12_port);
   M1_3_11 : MUX2_X1 port map( A => ML_int_3_11_port, B => ML_int_3_3_port, S 
                           => n10, Z => ML_int_4_11_port);
   M1_3_10 : MUX2_X1 port map( A => ML_int_3_10_port, B => ML_int_3_2_port, S 
                           => n10, Z => ML_int_4_10_port);
   M1_3_9 : MUX2_X1 port map( A => ML_int_3_9_port, B => ML_int_3_1_port, S => 
                           n10, Z => ML_int_4_9_port);
   M1_3_8 : MUX2_X1 port map( A => ML_int_3_8_port, B => ML_int_3_0_port, S => 
                           n10, Z => ML_int_4_8_port);
   M0_3_7 : MUX2_X1 port map( A => ML_int_3_7_port, B => ML_int_3_31_port, S =>
                           n10, Z => ML_int_4_7_port);
   M0_3_6 : MUX2_X1 port map( A => ML_int_3_6_port, B => ML_int_3_30_port, S =>
                           n10, Z => ML_int_4_6_port);
   M0_3_5 : MUX2_X1 port map( A => ML_int_3_5_port, B => ML_int_3_29_port, S =>
                           n10, Z => ML_int_4_5_port);
   M0_3_4 : MUX2_X1 port map( A => ML_int_3_4_port, B => ML_int_3_28_port, S =>
                           n10, Z => ML_int_4_4_port);
   M0_3_3 : MUX2_X1 port map( A => ML_int_3_3_port, B => ML_int_3_27_port, S =>
                           n10, Z => ML_int_4_3_port);
   M0_3_2 : MUX2_X1 port map( A => ML_int_3_2_port, B => ML_int_3_26_port, S =>
                           n10, Z => ML_int_4_2_port);
   M0_3_1 : MUX2_X1 port map( A => ML_int_3_1_port, B => ML_int_3_25_port, S =>
                           n10, Z => ML_int_4_1_port);
   M0_3_0 : MUX2_X1 port map( A => ML_int_3_0_port, B => ML_int_3_24_port, S =>
                           n10, Z => ML_int_4_0_port);
   M1_2_31 : MUX2_X1 port map( A => ML_int_2_31_port, B => ML_int_2_27_port, S 
                           => n9, Z => ML_int_3_31_port);
   M1_2_30 : MUX2_X1 port map( A => ML_int_2_30_port, B => ML_int_2_26_port, S 
                           => n9, Z => ML_int_3_30_port);
   M1_2_29 : MUX2_X1 port map( A => ML_int_2_29_port, B => ML_int_2_25_port, S 
                           => n9, Z => ML_int_3_29_port);
   M1_2_28 : MUX2_X1 port map( A => ML_int_2_28_port, B => ML_int_2_24_port, S 
                           => n9, Z => ML_int_3_28_port);
   M1_2_27 : MUX2_X1 port map( A => ML_int_2_27_port, B => ML_int_2_23_port, S 
                           => n9, Z => ML_int_3_27_port);
   M1_2_26 : MUX2_X1 port map( A => ML_int_2_26_port, B => ML_int_2_22_port, S 
                           => n9, Z => ML_int_3_26_port);
   M1_2_25 : MUX2_X1 port map( A => ML_int_2_25_port, B => ML_int_2_21_port, S 
                           => n9, Z => ML_int_3_25_port);
   M1_2_24 : MUX2_X1 port map( A => ML_int_2_24_port, B => ML_int_2_20_port, S 
                           => n9, Z => ML_int_3_24_port);
   M1_2_23 : MUX2_X1 port map( A => ML_int_2_23_port, B => ML_int_2_19_port, S 
                           => n8, Z => ML_int_3_23_port);
   M1_2_22 : MUX2_X1 port map( A => ML_int_2_22_port, B => ML_int_2_18_port, S 
                           => n8, Z => ML_int_3_22_port);
   M1_2_21 : MUX2_X1 port map( A => ML_int_2_21_port, B => ML_int_2_17_port, S 
                           => n8, Z => ML_int_3_21_port);
   M1_2_20 : MUX2_X1 port map( A => ML_int_2_20_port, B => ML_int_2_16_port, S 
                           => n8, Z => ML_int_3_20_port);
   M1_2_19 : MUX2_X1 port map( A => ML_int_2_19_port, B => ML_int_2_15_port, S 
                           => n8, Z => ML_int_3_19_port);
   M1_2_18 : MUX2_X1 port map( A => ML_int_2_18_port, B => ML_int_2_14_port, S 
                           => n8, Z => ML_int_3_18_port);
   M1_2_17 : MUX2_X1 port map( A => ML_int_2_17_port, B => ML_int_2_13_port, S 
                           => n8, Z => ML_int_3_17_port);
   M1_2_16 : MUX2_X1 port map( A => ML_int_2_16_port, B => ML_int_2_12_port, S 
                           => n8, Z => ML_int_3_16_port);
   M1_2_15 : MUX2_X1 port map( A => ML_int_2_15_port, B => ML_int_2_11_port, S 
                           => n8, Z => ML_int_3_15_port);
   M1_2_14 : MUX2_X1 port map( A => ML_int_2_14_port, B => ML_int_2_10_port, S 
                           => n8, Z => ML_int_3_14_port);
   M1_2_13 : MUX2_X1 port map( A => ML_int_2_13_port, B => ML_int_2_9_port, S 
                           => n8, Z => ML_int_3_13_port);
   M1_2_12 : MUX2_X1 port map( A => ML_int_2_12_port, B => ML_int_2_8_port, S 
                           => n8, Z => ML_int_3_12_port);
   M1_2_11 : MUX2_X1 port map( A => ML_int_2_11_port, B => ML_int_2_7_port, S 
                           => n7, Z => ML_int_3_11_port);
   M1_2_10 : MUX2_X1 port map( A => ML_int_2_10_port, B => ML_int_2_6_port, S 
                           => n7, Z => ML_int_3_10_port);
   M1_2_9 : MUX2_X1 port map( A => ML_int_2_9_port, B => ML_int_2_5_port, S => 
                           n7, Z => ML_int_3_9_port);
   M1_2_8 : MUX2_X1 port map( A => ML_int_2_8_port, B => ML_int_2_4_port, S => 
                           n7, Z => ML_int_3_8_port);
   M1_2_7 : MUX2_X1 port map( A => ML_int_2_7_port, B => ML_int_2_3_port, S => 
                           n7, Z => ML_int_3_7_port);
   M1_2_6 : MUX2_X1 port map( A => ML_int_2_6_port, B => ML_int_2_2_port, S => 
                           n7, Z => ML_int_3_6_port);
   M1_2_5 : MUX2_X1 port map( A => ML_int_2_5_port, B => ML_int_2_1_port, S => 
                           n7, Z => ML_int_3_5_port);
   M1_2_4 : MUX2_X1 port map( A => ML_int_2_4_port, B => ML_int_2_0_port, S => 
                           n7, Z => ML_int_3_4_port);
   M0_2_3 : MUX2_X1 port map( A => ML_int_2_3_port, B => ML_int_2_31_port, S =>
                           n7, Z => ML_int_3_3_port);
   M0_2_2 : MUX2_X1 port map( A => ML_int_2_2_port, B => ML_int_2_30_port, S =>
                           n7, Z => ML_int_3_2_port);
   M0_2_1 : MUX2_X1 port map( A => ML_int_2_1_port, B => ML_int_2_29_port, S =>
                           n7, Z => ML_int_3_1_port);
   M0_2_0 : MUX2_X1 port map( A => ML_int_2_0_port, B => ML_int_2_28_port, S =>
                           n7, Z => ML_int_3_0_port);
   M1_1_31 : MUX2_X1 port map( A => ML_int_1_31_port, B => ML_int_1_29_port, S 
                           => n6, Z => ML_int_2_31_port);
   M1_1_30 : MUX2_X1 port map( A => ML_int_1_30_port, B => ML_int_1_28_port, S 
                           => n6, Z => ML_int_2_30_port);
   M1_1_29 : MUX2_X1 port map( A => ML_int_1_29_port, B => ML_int_1_27_port, S 
                           => n6, Z => ML_int_2_29_port);
   M1_1_28 : MUX2_X1 port map( A => ML_int_1_28_port, B => ML_int_1_26_port, S 
                           => n6, Z => ML_int_2_28_port);
   M1_1_27 : MUX2_X1 port map( A => ML_int_1_27_port, B => ML_int_1_25_port, S 
                           => n6, Z => ML_int_2_27_port);
   M1_1_26 : MUX2_X1 port map( A => ML_int_1_26_port, B => ML_int_1_24_port, S 
                           => n6, Z => ML_int_2_26_port);
   M1_1_25 : MUX2_X1 port map( A => ML_int_1_25_port, B => ML_int_1_23_port, S 
                           => n6, Z => ML_int_2_25_port);
   M1_1_24 : MUX2_X1 port map( A => ML_int_1_24_port, B => ML_int_1_22_port, S 
                           => n6, Z => ML_int_2_24_port);
   M1_1_23 : MUX2_X1 port map( A => ML_int_1_23_port, B => ML_int_1_21_port, S 
                           => n5, Z => ML_int_2_23_port);
   M1_1_22 : MUX2_X1 port map( A => ML_int_1_22_port, B => ML_int_1_20_port, S 
                           => n5, Z => ML_int_2_22_port);
   M1_1_21 : MUX2_X1 port map( A => ML_int_1_21_port, B => ML_int_1_19_port, S 
                           => n5, Z => ML_int_2_21_port);
   M1_1_20 : MUX2_X1 port map( A => ML_int_1_20_port, B => ML_int_1_18_port, S 
                           => n5, Z => ML_int_2_20_port);
   M1_1_19 : MUX2_X1 port map( A => ML_int_1_19_port, B => ML_int_1_17_port, S 
                           => n5, Z => ML_int_2_19_port);
   M1_1_18 : MUX2_X1 port map( A => ML_int_1_18_port, B => ML_int_1_16_port, S 
                           => n5, Z => ML_int_2_18_port);
   M1_1_17 : MUX2_X1 port map( A => ML_int_1_17_port, B => ML_int_1_15_port, S 
                           => n5, Z => ML_int_2_17_port);
   M1_1_16 : MUX2_X1 port map( A => ML_int_1_16_port, B => ML_int_1_14_port, S 
                           => n5, Z => ML_int_2_16_port);
   M1_1_15 : MUX2_X1 port map( A => ML_int_1_15_port, B => ML_int_1_13_port, S 
                           => n5, Z => ML_int_2_15_port);
   M1_1_14 : MUX2_X1 port map( A => ML_int_1_14_port, B => ML_int_1_12_port, S 
                           => n5, Z => ML_int_2_14_port);
   M1_1_13 : MUX2_X1 port map( A => ML_int_1_13_port, B => ML_int_1_11_port, S 
                           => n5, Z => ML_int_2_13_port);
   M1_1_12 : MUX2_X1 port map( A => ML_int_1_12_port, B => ML_int_1_10_port, S 
                           => n5, Z => ML_int_2_12_port);
   M1_1_11 : MUX2_X1 port map( A => ML_int_1_11_port, B => ML_int_1_9_port, S 
                           => n4, Z => ML_int_2_11_port);
   M1_1_10 : MUX2_X1 port map( A => ML_int_1_10_port, B => ML_int_1_8_port, S 
                           => n4, Z => ML_int_2_10_port);
   M1_1_9 : MUX2_X1 port map( A => ML_int_1_9_port, B => ML_int_1_7_port, S => 
                           n4, Z => ML_int_2_9_port);
   M1_1_8 : MUX2_X1 port map( A => ML_int_1_8_port, B => ML_int_1_6_port, S => 
                           n4, Z => ML_int_2_8_port);
   M1_1_7 : MUX2_X1 port map( A => ML_int_1_7_port, B => ML_int_1_5_port, S => 
                           n4, Z => ML_int_2_7_port);
   M1_1_6 : MUX2_X1 port map( A => ML_int_1_6_port, B => ML_int_1_4_port, S => 
                           n4, Z => ML_int_2_6_port);
   M1_1_5 : MUX2_X1 port map( A => ML_int_1_5_port, B => ML_int_1_3_port, S => 
                           n4, Z => ML_int_2_5_port);
   M1_1_4 : MUX2_X1 port map( A => ML_int_1_4_port, B => ML_int_1_2_port, S => 
                           n4, Z => ML_int_2_4_port);
   M1_1_3 : MUX2_X1 port map( A => ML_int_1_3_port, B => ML_int_1_1_port, S => 
                           n4, Z => ML_int_2_3_port);
   M1_1_2 : MUX2_X1 port map( A => ML_int_1_2_port, B => ML_int_1_0_port, S => 
                           n4, Z => ML_int_2_2_port);
   M0_1_1 : MUX2_X1 port map( A => ML_int_1_1_port, B => ML_int_1_31_port, S =>
                           n4, Z => ML_int_2_1_port);
   M0_1_0 : MUX2_X1 port map( A => ML_int_1_0_port, B => ML_int_1_30_port, S =>
                           n4, Z => ML_int_2_0_port);
   M1_0_31 : MUX2_X1 port map( A => A(31), B => A(30), S => n3, Z => 
                           ML_int_1_31_port);
   M1_0_30 : MUX2_X1 port map( A => A(30), B => A(29), S => n3, Z => 
                           ML_int_1_30_port);
   M1_0_29 : MUX2_X1 port map( A => A(29), B => A(28), S => n3, Z => 
                           ML_int_1_29_port);
   M1_0_28 : MUX2_X1 port map( A => A(28), B => A(27), S => n3, Z => 
                           ML_int_1_28_port);
   M1_0_27 : MUX2_X1 port map( A => A(27), B => A(26), S => n3, Z => 
                           ML_int_1_27_port);
   M1_0_26 : MUX2_X1 port map( A => A(26), B => A(25), S => n3, Z => 
                           ML_int_1_26_port);
   M1_0_25 : MUX2_X1 port map( A => A(25), B => A(24), S => n3, Z => 
                           ML_int_1_25_port);
   M1_0_24 : MUX2_X1 port map( A => A(24), B => A(23), S => n3, Z => 
                           ML_int_1_24_port);
   M1_0_23 : MUX2_X1 port map( A => A(23), B => A(22), S => n2, Z => 
                           ML_int_1_23_port);
   M1_0_22 : MUX2_X1 port map( A => A(22), B => A(21), S => n2, Z => 
                           ML_int_1_22_port);
   M1_0_21 : MUX2_X1 port map( A => A(21), B => A(20), S => n2, Z => 
                           ML_int_1_21_port);
   M1_0_20 : MUX2_X1 port map( A => A(20), B => A(19), S => n2, Z => 
                           ML_int_1_20_port);
   M1_0_19 : MUX2_X1 port map( A => A(19), B => A(18), S => n2, Z => 
                           ML_int_1_19_port);
   M1_0_18 : MUX2_X1 port map( A => A(18), B => A(17), S => n2, Z => 
                           ML_int_1_18_port);
   M1_0_17 : MUX2_X1 port map( A => A(17), B => A(16), S => n2, Z => 
                           ML_int_1_17_port);
   M1_0_16 : MUX2_X1 port map( A => A(16), B => A(15), S => n2, Z => 
                           ML_int_1_16_port);
   M1_0_15 : MUX2_X1 port map( A => A(15), B => A(14), S => n2, Z => 
                           ML_int_1_15_port);
   M1_0_14 : MUX2_X1 port map( A => A(14), B => A(13), S => n2, Z => 
                           ML_int_1_14_port);
   M1_0_13 : MUX2_X1 port map( A => A(13), B => A(12), S => n2, Z => 
                           ML_int_1_13_port);
   M1_0_12 : MUX2_X1 port map( A => A(12), B => A(11), S => n2, Z => 
                           ML_int_1_12_port);
   M1_0_11 : MUX2_X1 port map( A => A(11), B => A(10), S => n1, Z => 
                           ML_int_1_11_port);
   M1_0_10 : MUX2_X1 port map( A => A(10), B => A(9), S => n1, Z => 
                           ML_int_1_10_port);
   M1_0_9 : MUX2_X1 port map( A => A(9), B => A(8), S => n1, Z => 
                           ML_int_1_9_port);
   M1_0_8 : MUX2_X1 port map( A => A(8), B => A(7), S => n1, Z => 
                           ML_int_1_8_port);
   M1_0_7 : MUX2_X1 port map( A => A(7), B => A(6), S => n1, Z => 
                           ML_int_1_7_port);
   M1_0_6 : MUX2_X1 port map( A => A(6), B => A(5), S => n1, Z => 
                           ML_int_1_6_port);
   M1_0_5 : MUX2_X1 port map( A => A(5), B => A(4), S => n1, Z => 
                           ML_int_1_5_port);
   M1_0_4 : MUX2_X1 port map( A => A(4), B => A(3), S => n1, Z => 
                           ML_int_1_4_port);
   M1_0_3 : MUX2_X1 port map( A => A(3), B => A(2), S => n1, Z => 
                           ML_int_1_3_port);
   M1_0_2 : MUX2_X1 port map( A => A(2), B => A(1), S => n1, Z => 
                           ML_int_1_2_port);
   M1_0_1 : MUX2_X1 port map( A => A(1), B => A(0), S => n1, Z => 
                           ML_int_1_1_port);
   M0_0_0 : MUX2_X1 port map( A => A(0), B => A(31), S => n1, Z => 
                           ML_int_1_0_port);
   U2 : BUF_X1 port map( A => SH(4), Z => n14);
   U3 : BUF_X1 port map( A => SH(4), Z => n13);
   U4 : BUF_X1 port map( A => SH(4), Z => n15);
   U5 : BUF_X1 port map( A => SH(1), Z => n5);
   U6 : BUF_X1 port map( A => SH(1), Z => n4);
   U7 : BUF_X1 port map( A => SH(2), Z => n8);
   U8 : BUF_X1 port map( A => SH(2), Z => n7);
   U9 : BUF_X1 port map( A => SH(0), Z => n2);
   U10 : BUF_X1 port map( A => SH(0), Z => n1);
   U11 : BUF_X1 port map( A => SH(3), Z => n11);
   U12 : BUF_X1 port map( A => SH(3), Z => n10);
   U13 : BUF_X1 port map( A => SH(1), Z => n6);
   U14 : BUF_X1 port map( A => SH(2), Z => n9);
   U15 : BUF_X1 port map( A => SH(0), Z => n3);
   U16 : BUF_X1 port map( A => SH(3), Z => n12);

end SYN_mx2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity SHIFTER_GENERIC_N32_DW_sra_0 is

   port( A : in std_logic_vector (31 downto 0);  SH : in std_logic_vector (4 
         downto 0);  SH_TC : in std_logic;  B : out std_logic_vector (31 downto
         0));

end SHIFTER_GENERIC_N32_DW_sra_0;

architecture SYN_mx2 of SHIFTER_GENERIC_N32_DW_sra_0 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component NOR2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal B_30_port, B_29_port, B_28_port, B_27_port, B_26_port, B_25_port, 
      B_24_port, B_23_port, B_22_port, B_21_port, B_20_port, B_19_port, 
      B_18_port, B_17_port, B_16_port, B_15_port, B_14_port, B_13_port, 
      B_12_port, B_11_port, B_10_port, B_9_port, B_8_port, B_7_port, B_6_port, 
      B_5_port, B_4_port, B_3_port, B_2_port, B_1_port, B_0_port, n1, n2, n3, 
      n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19,
      n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34
      , n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, 
      n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63
      , n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, 
      n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92
      , n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, 
      n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116, n117, 
      n118, n119, n120, n121, n122, n123, n124, n125, n126, n127, n128, n129, 
      n130, n131, n132, n133, n134, n135, n136, n137, n138, n139, n140, n141, 
      n142, n143, n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, 
      n154, n155, n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, 
      n166, n167, n168, n169, n170, n171, n172, n173, n174 : std_logic;

begin
   B <= ( A(31), B_30_port, B_29_port, B_28_port, B_27_port, B_26_port, 
      B_25_port, B_24_port, B_23_port, B_22_port, B_21_port, B_20_port, 
      B_19_port, B_18_port, B_17_port, B_16_port, B_15_port, B_14_port, 
      B_13_port, B_12_port, B_11_port, B_10_port, B_9_port, B_8_port, B_7_port,
      B_6_port, B_5_port, B_4_port, B_3_port, B_2_port, B_1_port, B_0_port );
   
   U2 : NOR2_X2 port map( A1 => n2, A2 => SH(0), ZN => n94);
   U3 : NOR2_X2 port map( A1 => SH(2), A2 => SH(3), ZN => n114);
   U4 : INV_X1 port map( A => n98, ZN => n59);
   U5 : INV_X1 port map( A => n95, ZN => n57);
   U6 : INV_X1 port map( A => n88, ZN => n54);
   U7 : INV_X1 port map( A => n4, ZN => n7);
   U8 : INV_X1 port map( A => n61, ZN => n55);
   U9 : INV_X1 port map( A => n97, ZN => n58);
   U10 : INV_X1 port map( A => n94, ZN => n56);
   U11 : NOR2_X2 port map( A1 => n1, A2 => n2, ZN => n95);
   U12 : NAND2_X1 port map( A1 => n1, A2 => n2, ZN => n98);
   U13 : AND2_X1 port map( A1 => n166, A2 => n3, ZN => n64);
   U14 : BUF_X1 port map( A => SH(4), Z => n4);
   U15 : BUF_X1 port map( A => SH(4), Z => n5);
   U16 : BUF_X1 port map( A => SH(4), Z => n6);
   U17 : INV_X1 port map( A => n121, ZN => n13);
   U18 : INV_X1 port map( A => n125, ZN => n11);
   U19 : INV_X1 port map( A => n126, ZN => n9);
   U20 : INV_X1 port map( A => n134, ZN => n15);
   U21 : INV_X1 port map( A => n138, ZN => n10);
   U22 : INV_X1 port map( A => n169, ZN => n8);
   U23 : INV_X1 port map( A => n137, ZN => n22);
   U24 : INV_X1 port map( A => n100, ZN => n16);
   U25 : INV_X1 port map( A => n141, ZN => n33);
   U26 : INV_X1 port map( A => n132, ZN => n34);
   U27 : INV_X1 port map( A => n149, ZN => n36);
   U28 : INV_X1 port map( A => n92, ZN => n38);
   U29 : INV_X1 port map( A => n104, ZN => n39);
   U30 : INV_X1 port map( A => n60, ZN => n41);
   U31 : INV_X1 port map( A => n68, ZN => n44);
   U32 : INV_X1 port map( A => n135, ZN => n14);
   U33 : INV_X1 port map( A => n77, ZN => n26);
   U34 : INV_X1 port map( A => n76, ZN => n30);
   U35 : INV_X1 port map( A => A(17), ZN => n32);
   U36 : INV_X1 port map( A => n168, ZN => n40);
   U37 : INV_X1 port map( A => A(12), ZN => n42);
   U38 : INV_X1 port map( A => n160, ZN => n35);
   U39 : INV_X1 port map( A => n148, ZN => n37);
   U40 : INV_X1 port map( A => A(21), ZN => n27);
   U41 : INV_X1 port map( A => A(23), ZN => n25);
   U42 : NAND2_X1 port map( A1 => n6, A2 => A(31), ZN => n100);
   U43 : INV_X1 port map( A => A(2), ZN => n53);
   U44 : INV_X1 port map( A => A(19), ZN => n29);
   U45 : INV_X1 port map( A => A(5), ZN => n50);
   U46 : INV_X1 port map( A => A(18), ZN => n31);
   U47 : INV_X1 port map( A => A(6), ZN => n49);
   U48 : INV_X1 port map( A => A(4), ZN => n51);
   U49 : INV_X1 port map( A => A(29), ZN => n18);
   U50 : INV_X1 port map( A => A(31), ZN => n12);
   U51 : INV_X1 port map( A => A(20), ZN => n28);
   U52 : INV_X1 port map( A => A(9), ZN => n46);
   U53 : INV_X1 port map( A => A(11), ZN => n43);
   U54 : INV_X1 port map( A => A(10), ZN => n45);
   U55 : INV_X1 port map( A => A(8), ZN => n47);
   U56 : INV_X1 port map( A => A(7), ZN => n48);
   U57 : INV_X1 port map( A => A(3), ZN => n52);
   U58 : INV_X1 port map( A => A(27), ZN => n20);
   U59 : INV_X1 port map( A => A(26), ZN => n21);
   U60 : INV_X1 port map( A => A(25), ZN => n23);
   U61 : INV_X1 port map( A => A(28), ZN => n19);
   U62 : INV_X1 port map( A => A(24), ZN => n24);
   U63 : INV_X1 port map( A => A(30), ZN => n17);
   U64 : INV_X1 port map( A => SH(0), ZN => n1);
   U65 : INV_X1 port map( A => SH(1), ZN => n2);
   U66 : INV_X1 port map( A => SH(2), ZN => n3);
   U67 : OAI221_X1 port map( B1 => n60, B2 => n61, C1 => n62, C2 => n7, A => 
                           n63, ZN => B_9_port);
   U68 : AOI222_X1 port map( A1 => n54, A2 => n34, B1 => n64, B2 => n65, C1 => 
                           n66, C2 => n67, ZN => n63);
   U69 : OAI221_X1 port map( B1 => n68, B2 => n61, C1 => n69, C2 => n7, A => 
                           n70, ZN => B_8_port);
   U70 : AOI222_X1 port map( A1 => n54, A2 => n36, B1 => n64, B2 => n71, C1 => 
                           n66, C2 => n72, ZN => n70);
   U71 : OAI221_X1 port map( B1 => n73, B2 => n61, C1 => n74, C2 => n7, A => 
                           n75, ZN => B_7_port);
   U72 : AOI222_X1 port map( A1 => n54, A2 => n38, B1 => n64, B2 => n76, C1 => 
                           n66, C2 => n77, ZN => n75);
   U73 : OAI221_X1 port map( B1 => n78, B2 => n61, C1 => n79, C2 => n7, A => 
                           n80, ZN => B_6_port);
   U74 : AOI222_X1 port map( A1 => n54, A2 => n39, B1 => n64, B2 => n33, C1 => 
                           n66, C2 => n81, ZN => n80);
   U75 : OAI221_X1 port map( B1 => n82, B2 => n61, C1 => n83, C2 => n7, A => 
                           n84, ZN => B_5_port);
   U76 : AOI222_X1 port map( A1 => n54, A2 => n41, B1 => n64, B2 => n34, C1 => 
                           n66, C2 => n65, ZN => n84);
   U77 : OAI221_X1 port map( B1 => n85, B2 => n61, C1 => n86, C2 => n7, A => 
                           n87, ZN => B_4_port);
   U78 : AOI222_X1 port map( A1 => n54, A2 => n44, B1 => n64, B2 => n36, C1 => 
                           n66, C2 => n71, ZN => n87);
   U79 : OAI221_X1 port map( B1 => n73, B2 => n88, C1 => n89, C2 => n7, A => 
                           n90, ZN => B_3_port);
   U80 : AOI222_X1 port map( A1 => n66, A2 => n76, B1 => n55, B2 => n91, C1 => 
                           n64, C2 => n38, ZN => n90);
   U81 : OAI221_X1 port map( B1 => n56, B2 => n50, C1 => n57, C2 => n49, A => 
                           n93, ZN => n91);
   U82 : AOI22_X1 port map( A1 => A(4), A2 => n58, B1 => A(3), B2 => n59, ZN =>
                           n93);
   U83 : AOI221_X1 port map( B1 => n94, B2 => A(9), C1 => n95, C2 => A(10), A 
                           => n96, ZN => n73);
   U84 : OAI22_X1 port map( A1 => n47, A2 => n97, B1 => n48, B2 => n98, ZN => 
                           n96);
   U85 : OAI21_X1 port map( B1 => n4, B2 => n99, A => n100, ZN => B_30_port);
   U86 : OAI221_X1 port map( B1 => n78, B2 => n88, C1 => n101, C2 => n7, A => 
                           n102, ZN => B_2_port);
   U87 : AOI222_X1 port map( A1 => n66, A2 => n33, B1 => n55, B2 => n103, C1 =>
                           n64, C2 => n39, ZN => n102);
   U88 : OAI221_X1 port map( B1 => n56, B2 => n51, C1 => n57, C2 => n50, A => 
                           n105, ZN => n103);
   U89 : AOI22_X1 port map( A1 => A(3), A2 => n58, B1 => A(2), B2 => n59, ZN =>
                           n105);
   U90 : AOI221_X1 port map( B1 => n94, B2 => A(8), C1 => n95, C2 => A(9), A =>
                           n106, ZN => n78);
   U91 : OAI22_X1 port map( A1 => n48, A2 => n97, B1 => n49, B2 => n98, ZN => 
                           n106);
   U92 : OAI21_X1 port map( B1 => n4, B2 => n107, A => n100, ZN => B_29_port);
   U93 : OAI21_X1 port map( B1 => n4, B2 => n108, A => n100, ZN => B_28_port);
   U94 : OAI21_X1 port map( B1 => n4, B2 => n109, A => n100, ZN => B_27_port);
   U95 : OAI21_X1 port map( B1 => n4, B2 => n110, A => n100, ZN => B_26_port);
   U96 : OAI21_X1 port map( B1 => n5, B2 => n62, A => n100, ZN => B_25_port);
   U97 : AOI221_X1 port map( B1 => n111, B2 => n112, C1 => n113, C2 => n114, A 
                           => n14, ZN => n62);
   U98 : OAI21_X1 port map( B1 => n5, B2 => n69, A => n100, ZN => B_24_port);
   U99 : AOI221_X1 port map( B1 => n115, B2 => n112, C1 => n116, C2 => n114, A 
                           => n14, ZN => n69);
   U100 : OAI21_X1 port map( B1 => n5, B2 => n74, A => n100, ZN => B_23_port);
   U101 : AOI221_X1 port map( B1 => n117, B2 => n112, C1 => n118, C2 => n114, A
                           => n14, ZN => n74);
   U102 : OAI21_X1 port map( B1 => n5, B2 => n79, A => n100, ZN => B_22_port);
   U103 : AOI221_X1 port map( B1 => n119, B2 => n112, C1 => n120, C2 => n114, A
                           => n13, ZN => n79);
   U104 : AOI21_X1 port map( B1 => n122, B2 => n123, A => n124, ZN => n121);
   U105 : OAI21_X1 port map( B1 => n5, B2 => n83, A => n100, ZN => B_21_port);
   U106 : AOI221_X1 port map( B1 => n113, B2 => n112, C1 => n67, C2 => n114, A 
                           => n11, ZN => n83);
   U107 : AOI21_X1 port map( B1 => n122, B2 => n111, A => n124, ZN => n125);
   U108 : OAI21_X1 port map( B1 => n5, B2 => n86, A => n100, ZN => B_20_port);
   U109 : AOI221_X1 port map( B1 => n116, B2 => n112, C1 => n72, C2 => n114, A 
                           => n9, ZN => n86);
   U110 : AOI21_X1 port map( B1 => n122, B2 => n115, A => n124, ZN => n126);
   U111 : OAI221_X1 port map( B1 => n82, B2 => n88, C1 => n127, C2 => n7, A => 
                           n128, ZN => B_1_port);
   U112 : AOI222_X1 port map( A1 => n66, A2 => n34, B1 => n55, B2 => n129, C1 
                           => n64, C2 => n41, ZN => n128);
   U113 : AOI221_X1 port map( B1 => n94, B2 => A(11), C1 => n95, C2 => A(12), A
                           => n130, ZN => n60);
   U114 : OAI22_X1 port map( A1 => n45, A2 => n97, B1 => n46, B2 => n98, ZN => 
                           n130);
   U115 : OAI221_X1 port map( B1 => n56, B2 => n52, C1 => n57, C2 => n51, A => 
                           n131, ZN => n129);
   U116 : AOI22_X1 port map( A1 => A(2), A2 => n58, B1 => A(1), B2 => n59, ZN 
                           => n131);
   U117 : AOI221_X1 port map( B1 => n94, B2 => A(7), C1 => n95, C2 => A(8), A 
                           => n133, ZN => n82);
   U118 : OAI22_X1 port map( A1 => n49, A2 => n97, B1 => n50, B2 => n98, ZN => 
                           n133);
   U119 : OAI21_X1 port map( B1 => n5, B2 => n89, A => n100, ZN => B_19_port);
   U120 : AOI221_X1 port map( B1 => n118, B2 => n112, C1 => n77, C2 => n114, A 
                           => n15, ZN => n89);
   U121 : AOI21_X1 port map( B1 => n122, B2 => n117, A => n124, ZN => n134);
   U122 : NOR2_X1 port map( A1 => n135, A2 => n3, ZN => n124);
   U123 : OAI21_X1 port map( B1 => n6, B2 => n101, A => n100, ZN => B_18_port);
   U124 : AOI221_X1 port map( B1 => n123, B2 => n136, C1 => n119, C2 => n122, A
                           => n22, ZN => n101);
   U125 : AOI22_X1 port map( A1 => n112, A2 => n120, B1 => n114, B2 => n81, ZN 
                           => n137);
   U126 : OAI21_X1 port map( B1 => n6, B2 => n127, A => n100, ZN => B_17_port);
   U127 : AOI221_X1 port map( B1 => n67, B2 => n112, C1 => n65, C2 => n114, A 
                           => n10, ZN => n127);
   U128 : AOI22_X1 port map( A1 => n136, A2 => n111, B1 => n122, B2 => n113, ZN
                           => n138);
   U129 : OAI21_X1 port map( B1 => n6, B2 => n139, A => n100, ZN => B_16_port);
   U130 : OAI221_X1 port map( B1 => n26, B2 => n88, C1 => n30, C2 => n61, A => 
                           n140, ZN => B_15_port);
   U131 : AOI221_X1 port map( B1 => n66, B2 => n117, C1 => n64, C2 => n118, A 
                           => n16, ZN => n140);
   U132 : OAI221_X1 port map( B1 => n141, B2 => n61, C1 => n99, C2 => n7, A => 
                           n142, ZN => B_14_port);
   U133 : AOI222_X1 port map( A1 => n54, A2 => n81, B1 => n64, B2 => n120, C1 
                           => n66, C2 => n119, ZN => n142);
   U134 : AOI21_X1 port map( B1 => n123, B2 => n114, A => n143, ZN => n99);
   U135 : OAI221_X1 port map( B1 => n132, B2 => n61, C1 => n107, C2 => n7, A =>
                           n144, ZN => B_13_port);
   U136 : AOI222_X1 port map( A1 => n54, A2 => n65, B1 => n64, B2 => n67, C1 =>
                           n66, C2 => n113, ZN => n144);
   U137 : OAI221_X1 port map( B1 => n56, B2 => n20, C1 => n57, C2 => n19, A => 
                           n145, ZN => n113);
   U138 : AOI22_X1 port map( A1 => A(26), A2 => n58, B1 => A(25), B2 => n59, ZN
                           => n145);
   U139 : OAI221_X1 port map( B1 => n56, B2 => n25, C1 => n57, C2 => n24, A => 
                           n146, ZN => n67);
   U140 : AOI22_X1 port map( A1 => A(22), A2 => n58, B1 => A(21), B2 => n59, ZN
                           => n146);
   U141 : OAI221_X1 port map( B1 => n56, B2 => n29, C1 => n57, C2 => n28, A => 
                           n147, ZN => n65);
   U142 : AOI22_X1 port map( A1 => A(18), A2 => n58, B1 => A(17), B2 => n59, ZN
                           => n147);
   U143 : AOI21_X1 port map( B1 => n111, B2 => n114, A => n143, ZN => n107);
   U144 : OAI222_X1 port map( A1 => n98, A2 => n18, B1 => n97, B2 => n17, C1 =>
                           n2, C2 => n12, ZN => n111);
   U145 : AOI221_X1 port map( B1 => n94, B2 => A(15), C1 => n95, C2 => A(16), A
                           => n37, ZN => n132);
   U146 : AOI22_X1 port map( A1 => A(14), A2 => n58, B1 => A(13), B2 => n59, ZN
                           => n148);
   U147 : OAI221_X1 port map( B1 => n149, B2 => n61, C1 => n108, C2 => n7, A =>
                           n150, ZN => B_12_port);
   U148 : AOI222_X1 port map( A1 => n54, A2 => n71, B1 => n64, B2 => n72, C1 =>
                           n66, C2 => n116, ZN => n150);
   U149 : AOI21_X1 port map( B1 => n115, B2 => n114, A => n143, ZN => n108);
   U150 : OAI221_X1 port map( B1 => n92, B2 => n61, C1 => n109, C2 => n7, A => 
                           n151, ZN => B_11_port);
   U151 : AOI222_X1 port map( A1 => n54, A2 => n76, B1 => n64, B2 => n77, C1 =>
                           n66, C2 => n118, ZN => n151);
   U152 : OAI221_X1 port map( B1 => n56, B2 => n23, C1 => n57, C2 => n21, A => 
                           n152, ZN => n118);
   U153 : AOI22_X1 port map( A1 => A(24), A2 => n58, B1 => A(23), B2 => n59, ZN
                           => n152);
   U154 : OAI221_X1 port map( B1 => n28, B2 => n97, C1 => n29, C2 => n98, A => 
                           n153, ZN => n77);
   U155 : AOI22_X1 port map( A1 => A(21), A2 => n94, B1 => A(22), B2 => n95, ZN
                           => n153);
   U156 : OAI221_X1 port map( B1 => n56, B2 => n32, C1 => n57, C2 => n31, A => 
                           n154, ZN => n76);
   U157 : AOI22_X1 port map( A1 => A(16), A2 => n58, B1 => A(15), B2 => n59, ZN
                           => n154);
   U158 : AOI21_X1 port map( B1 => n117, B2 => n114, A => n143, ZN => n109);
   U159 : OAI21_X1 port map( B1 => n3, B2 => n12, A => n135, ZN => n143);
   U160 : OAI221_X1 port map( B1 => n56, B2 => n18, C1 => n57, C2 => n17, A => 
                           n155, ZN => n117);
   U161 : AOI22_X1 port map( A1 => A(28), A2 => n58, B1 => A(27), B2 => n59, ZN
                           => n155);
   U162 : AOI221_X1 port map( B1 => n94, B2 => A(13), C1 => n95, C2 => A(14), A
                           => n156, ZN => n92);
   U163 : OAI22_X1 port map( A1 => n42, A2 => n97, B1 => n43, B2 => n98, ZN => 
                           n156);
   U164 : OAI221_X1 port map( B1 => n104, B2 => n61, C1 => n110, C2 => n7, A =>
                           n157, ZN => B_10_port);
   U165 : AOI222_X1 port map( A1 => n54, A2 => n33, B1 => n64, B2 => n81, C1 =>
                           n66, C2 => n120, ZN => n157);
   U166 : OAI221_X1 port map( B1 => n56, B2 => n24, C1 => n57, C2 => n23, A => 
                           n158, ZN => n120);
   U167 : AOI22_X1 port map( A1 => A(23), A2 => n58, B1 => A(22), B2 => n59, ZN
                           => n158);
   U168 : OAI221_X1 port map( B1 => n29, B2 => n97, C1 => n31, C2 => n98, A => 
                           n159, ZN => n81);
   U169 : AOI22_X1 port map( A1 => A(20), A2 => n94, B1 => A(21), B2 => n95, ZN
                           => n159);
   U170 : AOI221_X1 port map( B1 => n94, B2 => A(16), C1 => n95, C2 => A(17), A
                           => n35, ZN => n141);
   U171 : AOI22_X1 port map( A1 => A(15), A2 => n58, B1 => A(14), B2 => n59, ZN
                           => n160);
   U172 : AOI221_X1 port map( B1 => n123, B2 => n112, C1 => n119, C2 => n114, A
                           => n14, ZN => n110);
   U173 : NAND2_X1 port map( A1 => A(31), A2 => SH(3), ZN => n135);
   U174 : OAI221_X1 port map( B1 => n56, B2 => n19, C1 => n57, C2 => n18, A => 
                           n161, ZN => n119);
   U175 : AOI22_X1 port map( A1 => A(27), A2 => n58, B1 => A(26), B2 => n59, ZN
                           => n161);
   U176 : MUX2_X1 port map( A => A(30), B => A(31), S => n98, Z => n123);
   U177 : AOI221_X1 port map( B1 => n94, B2 => A(12), C1 => n95, C2 => A(13), A
                           => n162, ZN => n104);
   U178 : OAI22_X1 port map( A1 => n43, A2 => n97, B1 => n45, B2 => n98, ZN => 
                           n162);
   U179 : OAI221_X1 port map( B1 => n85, B2 => n88, C1 => n139, C2 => n7, A => 
                           n163, ZN => B_0_port);
   U180 : AOI222_X1 port map( A1 => n66, A2 => n36, B1 => n55, B2 => n164, C1 
                           => n64, C2 => n44, ZN => n163);
   U181 : AOI221_X1 port map( B1 => n94, B2 => A(10), C1 => n95, C2 => A(11), A
                           => n165, ZN => n68);
   U182 : OAI22_X1 port map( A1 => n46, A2 => n97, B1 => n47, B2 => n98, ZN => 
                           n165);
   U183 : OAI221_X1 port map( B1 => n56, B2 => n53, C1 => n57, C2 => n52, A => 
                           n167, ZN => n164);
   U184 : AOI22_X1 port map( A1 => A(1), A2 => n58, B1 => A(0), B2 => n59, ZN 
                           => n167);
   U185 : NAND2_X1 port map( A1 => n114, A2 => n7, ZN => n61);
   U186 : AOI221_X1 port map( B1 => n94, B2 => A(14), C1 => n95, C2 => A(15), A
                           => n40, ZN => n149);
   U187 : AOI22_X1 port map( A1 => A(13), A2 => n58, B1 => A(12), B2 => n59, ZN
                           => n168);
   U188 : AND2_X1 port map( A1 => SH(2), A2 => n166, ZN => n66);
   U189 : AND2_X1 port map( A1 => SH(3), A2 => n7, ZN => n166);
   U190 : AOI221_X1 port map( B1 => n72, B2 => n112, C1 => n71, C2 => n114, A 
                           => n8, ZN => n139);
   U191 : AOI22_X1 port map( A1 => n136, A2 => n115, B1 => n122, B2 => n116, ZN
                           => n169);
   U192 : OAI221_X1 port map( B1 => n56, B2 => n21, C1 => n57, C2 => n20, A => 
                           n170, ZN => n116);
   U193 : AOI22_X1 port map( A1 => A(25), A2 => n58, B1 => A(24), B2 => n59, ZN
                           => n170);
   U194 : AND2_X1 port map( A1 => SH(3), A2 => n3, ZN => n122);
   U195 : OAI221_X1 port map( B1 => n56, B2 => n17, C1 => n57, C2 => n12, A => 
                           n171, ZN => n115);
   U196 : AOI22_X1 port map( A1 => A(29), A2 => n58, B1 => A(28), B2 => n59, ZN
                           => n171);
   U197 : AND2_X1 port map( A1 => SH(2), A2 => SH(3), ZN => n136);
   U198 : OAI221_X1 port map( B1 => n56, B2 => n31, C1 => n29, C2 => n57, A => 
                           n172, ZN => n71);
   U199 : AOI22_X1 port map( A1 => A(17), A2 => n58, B1 => A(16), B2 => n59, ZN
                           => n172);
   U200 : OAI221_X1 port map( B1 => n97, B2 => n27, C1 => n28, C2 => n98, A => 
                           n173, ZN => n72);
   U201 : AOI22_X1 port map( A1 => A(22), A2 => n94, B1 => A(23), B2 => n95, ZN
                           => n173);
   U202 : NAND2_X1 port map( A1 => n112, A2 => n7, ZN => n88);
   U203 : NOR2_X1 port map( A1 => n3, A2 => SH(3), ZN => n112);
   U204 : AOI221_X1 port map( B1 => n94, B2 => A(6), C1 => n95, C2 => A(7), A 
                           => n174, ZN => n85);
   U205 : OAI22_X1 port map( A1 => n50, A2 => n97, B1 => n51, B2 => n98, ZN => 
                           n174);
   U206 : NAND2_X1 port map( A1 => SH(0), A2 => n2, ZN => n97);

end SYN_mx2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity SHIFTER_GENERIC_N32_DW_rash_0 is

   port( A : in std_logic_vector (31 downto 0);  DATA_TC : in std_logic;  SH : 
         in std_logic_vector (4 downto 0);  SH_TC : in std_logic;  B : out 
         std_logic_vector (31 downto 0));

end SHIFTER_GENERIC_N32_DW_rash_0;

architecture SYN_mx2 of SHIFTER_GENERIC_N32_DW_rash_0 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n12, n13, n14, n15, n16, n17
      , n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, 
      n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46
      , n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, 
      n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75
      , n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, 
      n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103,
      n104, n105, n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, 
      n116, n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, n127, 
      n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, n138, n139, 
      n140, n141, n142, n143, n144, n145, n146, n147, n148, n149, n150, n151, 
      n152, n153, n154, n155, n156, n157, n158, n159, n160, n161, n162, n163, 
      n164, n165, n166, n167, n168 : std_logic;

begin
   
   U3 : INV_X1 port map( A => n62, ZN => n55);
   U4 : INV_X1 port map( A => n143, ZN => n56);
   U5 : INV_X1 port map( A => n8, ZN => n9);
   U6 : INV_X1 port map( A => n92, ZN => n54);
   U7 : INV_X1 port map( A => n97, ZN => n60);
   U8 : INV_X1 port map( A => n101, ZN => n57);
   U9 : INV_X1 port map( A => n100, ZN => n58);
   U10 : INV_X1 port map( A => n98, ZN => n59);
   U11 : AND2_X1 port map( A1 => n160, A2 => n4, ZN => n66);
   U12 : BUF_X1 port map( A => SH(4), Z => n8);
   U13 : BUF_X1 port map( A => SH(4), Z => n6);
   U14 : BUF_X1 port map( A => SH(4), Z => n7);
   U15 : BUF_X1 port map( A => n98, Z => n1);
   U16 : BUF_X1 port map( A => n98, Z => n2);
   U17 : INV_X1 port map( A => n128, ZN => n14);
   U18 : NOR2_X2 port map( A1 => n3, A2 => SH(1), ZN => n100);
   U19 : INV_X1 port map( A => n129, ZN => n13);
   U20 : INV_X1 port map( A => n131, ZN => n15);
   U21 : INV_X1 port map( A => n163, ZN => n10);
   U22 : INV_X1 port map( A => n142, ZN => n12);
   U23 : INV_X1 port map( A => n141, ZN => B(12));
   U24 : INV_X1 port map( A => n61, ZN => n41);
   U25 : INV_X1 port map( A => n79, ZN => n31);
   U26 : INV_X1 port map( A => n108, ZN => n40);
   U27 : INV_X1 port map( A => n70, ZN => n44);
   U28 : INV_X1 port map( A => n96, ZN => n38);
   U29 : INV_X1 port map( A => n84, ZN => n33);
   U30 : INV_X1 port map( A => n65, ZN => n35);
   U31 : INV_X1 port map( A => n85, ZN => n26);
   U32 : INV_X1 port map( A => n67, ZN => n28);
   U33 : INV_X1 port map( A => n80, ZN => n25);
   U34 : INV_X1 port map( A => A(14), ZN => n39);
   U35 : INV_X1 port map( A => A(23), ZN => n24);
   U36 : INV_X1 port map( A => A(12), ZN => n42);
   U37 : INV_X1 port map( A => A(2), ZN => n53);
   U38 : INV_X1 port map( A => A(31), ZN => n16);
   U39 : INV_X1 port map( A => A(20), ZN => n29);
   U40 : INV_X1 port map( A => A(5), ZN => n50);
   U41 : INV_X1 port map( A => A(30), ZN => n17);
   U42 : INV_X1 port map( A => A(6), ZN => n49);
   U43 : INV_X1 port map( A => A(4), ZN => n51);
   U44 : INV_X1 port map( A => A(29), ZN => n18);
   U45 : INV_X1 port map( A => A(19), ZN => n30);
   U46 : INV_X1 port map( A => A(17), ZN => n34);
   U47 : INV_X1 port map( A => A(21), ZN => n27);
   U48 : INV_X1 port map( A => A(9), ZN => n46);
   U49 : INV_X1 port map( A => A(11), ZN => n43);
   U50 : INV_X1 port map( A => A(10), ZN => n45);
   U51 : INV_X1 port map( A => A(8), ZN => n47);
   U52 : INV_X1 port map( A => A(7), ZN => n48);
   U53 : INV_X1 port map( A => A(16), ZN => n36);
   U54 : INV_X1 port map( A => A(15), ZN => n37);
   U55 : INV_X1 port map( A => A(3), ZN => n52);
   U56 : INV_X1 port map( A => A(26), ZN => n21);
   U57 : INV_X1 port map( A => A(27), ZN => n20);
   U58 : INV_X1 port map( A => A(28), ZN => n19);
   U59 : INV_X1 port map( A => A(25), ZN => n22);
   U60 : INV_X1 port map( A => A(24), ZN => n23);
   U61 : INV_X1 port map( A => A(18), ZN => n32);
   U62 : NOR2_X2 port map( A1 => SH(0), A2 => SH(1), ZN => n101);
   U63 : INV_X1 port map( A => SH(0), ZN => n3);
   U64 : INV_X1 port map( A => SH(2), ZN => n4);
   U65 : INV_X1 port map( A => SH(3), ZN => n5);
   U66 : OAI221_X1 port map( B1 => n61, B2 => n62, C1 => n63, C2 => n9, A => 
                           n64, ZN => B(9));
   U67 : AOI222_X1 port map( A1 => n54, A2 => n65, B1 => n66, B2 => n67, C1 => 
                           n68, C2 => n69, ZN => n64);
   U68 : OAI221_X1 port map( B1 => n70, B2 => n62, C1 => n71, C2 => n9, A => 
                           n72, ZN => B(8));
   U69 : AOI222_X1 port map( A1 => n54, A2 => n73, B1 => n66, B2 => n74, C1 => 
                           n68, C2 => n75, ZN => n72);
   U70 : OAI221_X1 port map( B1 => n76, B2 => n62, C1 => n77, C2 => n9, A => 
                           n78, ZN => B(7));
   U71 : AOI222_X1 port map( A1 => n54, A2 => n38, B1 => n66, B2 => n79, C1 => 
                           n68, C2 => n80, ZN => n78);
   U72 : OAI221_X1 port map( B1 => n81, B2 => n62, C1 => n82, C2 => n9, A => 
                           n83, ZN => B(6));
   U73 : AOI222_X1 port map( A1 => n54, A2 => n40, B1 => n66, B2 => n84, C1 => 
                           n68, C2 => n85, ZN => n83);
   U74 : OAI221_X1 port map( B1 => n86, B2 => n62, C1 => n87, C2 => n9, A => 
                           n88, ZN => B(5));
   U75 : AOI222_X1 port map( A1 => n54, A2 => n41, B1 => n66, B2 => n65, C1 => 
                           n68, C2 => n67, ZN => n88);
   U76 : OAI221_X1 port map( B1 => n89, B2 => n62, C1 => n90, C2 => n9, A => 
                           n91, ZN => B(4));
   U77 : AOI222_X1 port map( A1 => n54, A2 => n44, B1 => n66, B2 => n73, C1 => 
                           n68, C2 => n74, ZN => n91);
   U78 : OAI221_X1 port map( B1 => n76, B2 => n92, C1 => n93, C2 => n9, A => 
                           n94, ZN => B(3));
   U79 : AOI222_X1 port map( A1 => n68, A2 => n79, B1 => n55, B2 => n95, C1 => 
                           n66, C2 => n38, ZN => n94);
   U80 : OAI221_X1 port map( B1 => n97, B2 => n49, C1 => n1, C2 => n50, A => 
                           n99, ZN => n95);
   U81 : AOI22_X1 port map( A1 => A(4), A2 => n100, B1 => A(3), B2 => n101, ZN 
                           => n99);
   U82 : AOI221_X1 port map( B1 => n60, B2 => A(10), C1 => n59, C2 => A(9), A 
                           => n102, ZN => n76);
   U83 : OAI22_X1 port map( A1 => n47, A2 => n58, B1 => n48, B2 => n57, ZN => 
                           n102);
   U84 : AND2_X1 port map( A1 => n55, A2 => n103, ZN => B(31));
   U85 : AND2_X1 port map( A1 => n104, A2 => n55, ZN => B(30));
   U86 : OAI221_X1 port map( B1 => n81, B2 => n92, C1 => n105, C2 => n9, A => 
                           n106, ZN => B(2));
   U87 : AOI222_X1 port map( A1 => n68, A2 => n84, B1 => n55, B2 => n107, C1 =>
                           n66, C2 => n40, ZN => n106);
   U88 : OAI221_X1 port map( B1 => n97, B2 => n50, C1 => n2, C2 => n51, A => 
                           n109, ZN => n107);
   U89 : AOI22_X1 port map( A1 => A(3), A2 => n100, B1 => A(2), B2 => n101, ZN 
                           => n109);
   U90 : AOI221_X1 port map( B1 => n60, B2 => A(9), C1 => n59, C2 => A(8), A =>
                           n110, ZN => n81);
   U91 : OAI22_X1 port map( A1 => n48, A2 => n58, B1 => n49, B2 => n57, ZN => 
                           n110);
   U92 : AND2_X1 port map( A1 => n111, A2 => n55, ZN => B(29));
   U93 : AND2_X1 port map( A1 => n112, A2 => n55, ZN => B(28));
   U94 : NOR3_X1 port map( A1 => n14, A2 => n8, A3 => SH(3), ZN => B(27));
   U95 : NOR2_X1 port map( A1 => n6, A2 => n113, ZN => B(26));
   U96 : NOR2_X1 port map( A1 => n6, A2 => n63, ZN => B(25));
   U97 : AOI22_X1 port map( A1 => n114, A2 => n56, B1 => n111, B2 => n115, ZN 
                           => n63);
   U98 : NOR2_X1 port map( A1 => n6, A2 => n71, ZN => B(24));
   U99 : AOI22_X1 port map( A1 => n116, A2 => n56, B1 => n112, B2 => n115, ZN 
                           => n71);
   U100 : NOR2_X1 port map( A1 => n6, A2 => n77, ZN => B(23));
   U101 : AOI222_X1 port map( A1 => n117, A2 => n115, B1 => n103, B2 => n118, 
                           C1 => n119, C2 => n56, ZN => n77);
   U102 : NOR2_X1 port map( A1 => n6, A2 => n82, ZN => B(22));
   U103 : AOI222_X1 port map( A1 => n120, A2 => n115, B1 => n104, B2 => n118, 
                           C1 => n121, C2 => n56, ZN => n82);
   U104 : NOR2_X1 port map( A1 => n7, A2 => n87, ZN => B(21));
   U105 : AOI222_X1 port map( A1 => n114, A2 => n115, B1 => n111, B2 => n118, 
                           C1 => n69, C2 => n56, ZN => n87);
   U106 : NOR2_X1 port map( A1 => n7, A2 => n90, ZN => B(20));
   U107 : AOI222_X1 port map( A1 => n116, A2 => n115, B1 => n112, B2 => n118, 
                           C1 => n75, C2 => n56, ZN => n90);
   U108 : OAI221_X1 port map( B1 => n86, B2 => n92, C1 => n122, C2 => n9, A => 
                           n123, ZN => B(1));
   U109 : AOI222_X1 port map( A1 => n68, A2 => n65, B1 => n55, B2 => n124, C1 
                           => n66, C2 => n41, ZN => n123);
   U110 : AOI221_X1 port map( B1 => n60, B2 => A(12), C1 => n59, C2 => A(11), A
                           => n125, ZN => n61);
   U111 : OAI22_X1 port map( A1 => n45, A2 => n58, B1 => n46, B2 => n57, ZN => 
                           n125);
   U112 : OAI221_X1 port map( B1 => n97, B2 => n51, C1 => n2, C2 => n52, A => 
                           n126, ZN => n124);
   U113 : AOI22_X1 port map( A1 => A(2), A2 => n100, B1 => A(1), B2 => n101, ZN
                           => n126);
   U114 : AOI221_X1 port map( B1 => n60, B2 => A(8), C1 => n59, C2 => A(7), A 
                           => n127, ZN => n86);
   U115 : OAI22_X1 port map( A1 => n49, A2 => n58, B1 => n50, B2 => n57, ZN => 
                           n127);
   U116 : NOR2_X1 port map( A1 => n7, A2 => n93, ZN => B(19));
   U117 : AOI222_X1 port map( A1 => n80, A2 => n56, B1 => n119, B2 => n115, C1 
                           => n128, C2 => SH(3), ZN => n93);
   U118 : NOR2_X1 port map( A1 => n7, A2 => n105, ZN => B(18));
   U119 : AOI221_X1 port map( B1 => n121, B2 => n115, C1 => n85, C2 => n56, A 
                           => n13, ZN => n105);
   U120 : AOI22_X1 port map( A1 => n130, A2 => n104, B1 => n118, B2 => n120, ZN
                           => n129);
   U121 : NOR2_X1 port map( A1 => n7, A2 => n122, ZN => B(17));
   U122 : AOI221_X1 port map( B1 => n69, B2 => n115, C1 => n67, C2 => n56, A =>
                           n15, ZN => n122);
   U123 : AOI22_X1 port map( A1 => n130, A2 => n111, B1 => n118, B2 => n114, ZN
                           => n131);
   U124 : NOR2_X1 port map( A1 => n8, A2 => n132, ZN => B(16));
   U125 : OAI221_X1 port map( B1 => n25, B2 => n92, C1 => n31, C2 => n62, A => 
                           n133, ZN => B(15));
   U126 : AOI222_X1 port map( A1 => n68, A2 => n117, B1 => n134, B2 => n103, C1
                           => n66, C2 => n119, ZN => n133);
   U127 : OAI221_X1 port map( B1 => n26, B2 => n92, C1 => n33, C2 => n62, A => 
                           n135, ZN => B(14));
   U128 : AOI222_X1 port map( A1 => n68, A2 => n120, B1 => n134, B2 => n104, C1
                           => n66, C2 => n121, ZN => n135);
   U129 : OAI221_X1 port map( B1 => n28, B2 => n92, C1 => n35, C2 => n62, A => 
                           n136, ZN => B(13));
   U130 : AOI222_X1 port map( A1 => n68, A2 => n114, B1 => n134, B2 => n111, C1
                           => n66, C2 => n69, ZN => n136);
   U131 : OAI221_X1 port map( B1 => n97, B2 => n23, C1 => n1, C2 => n24, A => 
                           n137, ZN => n69);
   U132 : AOI22_X1 port map( A1 => A(22), A2 => n100, B1 => A(21), B2 => n101, 
                           ZN => n137);
   U133 : OAI222_X1 port map( A1 => n58, A2 => n17, B1 => n1, B2 => n16, C1 => 
                           n57, C2 => n18, ZN => n111);
   U134 : OAI221_X1 port map( B1 => n97, B2 => n19, C1 => n1, C2 => n20, A => 
                           n138, ZN => n114);
   U135 : AOI22_X1 port map( A1 => A(26), A2 => n100, B1 => A(25), B2 => n101, 
                           ZN => n138);
   U136 : OAI221_X1 port map( B1 => n97, B2 => n36, C1 => n2, C2 => n37, A => 
                           n139, ZN => n65);
   U137 : AOI22_X1 port map( A1 => A(14), A2 => n100, B1 => A(13), B2 => n101, 
                           ZN => n139);
   U138 : OAI221_X1 port map( B1 => n97, B2 => n29, C1 => n2, C2 => n30, A => 
                           n140, ZN => n67);
   U139 : AOI22_X1 port map( A1 => A(18), A2 => n100, B1 => A(17), B2 => n101, 
                           ZN => n140);
   U140 : AOI221_X1 port map( B1 => n74, B2 => n54, C1 => n73, C2 => n55, A => 
                           n12, ZN => n141);
   U141 : AOI222_X1 port map( A1 => n68, A2 => n116, B1 => n134, B2 => n112, C1
                           => n66, C2 => n75, ZN => n142);
   U142 : NOR2_X1 port map( A1 => n9, A2 => n143, ZN => n134);
   U143 : OAI221_X1 port map( B1 => n31, B2 => n92, C1 => n96, C2 => n62, A => 
                           n144, ZN => B(11));
   U144 : AOI221_X1 port map( B1 => n68, B2 => n119, C1 => n66, C2 => n80, A =>
                           n145, ZN => n144);
   U145 : NOR3_X1 port map( A1 => n9, A2 => SH(3), A3 => n14, ZN => n145);
   U146 : MUX2_X1 port map( A => n117, B => n103, S => SH(2), Z => n128);
   U147 : NOR2_X1 port map( A1 => n16, A2 => n57, ZN => n103);
   U148 : OAI221_X1 port map( B1 => n97, B2 => n17, C1 => n1, C2 => n18, A => 
                           n146, ZN => n117);
   U149 : AOI22_X1 port map( A1 => A(28), A2 => n100, B1 => A(27), B2 => n101, 
                           ZN => n146);
   U150 : OAI221_X1 port map( B1 => n29, B2 => n58, C1 => n30, C2 => n57, A => 
                           n147, ZN => n80);
   U151 : AOI22_X1 port map( A1 => A(22), A2 => n60, B1 => A(21), B2 => n59, ZN
                           => n147);
   U152 : OAI221_X1 port map( B1 => n97, B2 => n21, C1 => n1, C2 => n22, A => 
                           n148, ZN => n119);
   U153 : AOI22_X1 port map( A1 => A(24), A2 => n100, B1 => A(23), B2 => n101, 
                           ZN => n148);
   U154 : AOI221_X1 port map( B1 => n60, B2 => A(14), C1 => n59, C2 => A(13), A
                           => n149, ZN => n96);
   U155 : OAI22_X1 port map( A1 => n42, A2 => n58, B1 => n43, B2 => n57, ZN => 
                           n149);
   U156 : OAI221_X1 port map( B1 => n97, B2 => n32, C1 => n2, C2 => n34, A => 
                           n150, ZN => n79);
   U157 : AOI22_X1 port map( A1 => A(16), A2 => n100, B1 => A(15), B2 => n101, 
                           ZN => n150);
   U158 : OAI221_X1 port map( B1 => n108, B2 => n62, C1 => n113, C2 => n9, A =>
                           n151, ZN => B(10));
   U159 : AOI222_X1 port map( A1 => n54, A2 => n84, B1 => n66, B2 => n85, C1 =>
                           n68, C2 => n121, ZN => n151);
   U160 : OAI221_X1 port map( B1 => n97, B2 => n22, C1 => n2, C2 => n23, A => 
                           n152, ZN => n121);
   U161 : AOI22_X1 port map( A1 => A(23), A2 => n100, B1 => A(22), B2 => n101, 
                           ZN => n152);
   U162 : OAI221_X1 port map( B1 => n97, B2 => n27, C1 => n29, C2 => n2, A => 
                           n153, ZN => n85);
   U163 : AOI22_X1 port map( A1 => n100, A2 => A(19), B1 => n101, B2 => A(18), 
                           ZN => n153);
   U164 : OAI221_X1 port map( B1 => n97, B2 => n34, C1 => n1, C2 => n36, A => 
                           n154, ZN => n84);
   U165 : AOI22_X1 port map( A1 => A(15), A2 => n100, B1 => A(14), B2 => n101, 
                           ZN => n154);
   U166 : AOI22_X1 port map( A1 => n120, A2 => n56, B1 => n104, B2 => n115, ZN 
                           => n113);
   U167 : OAI22_X1 port map( A1 => n57, A2 => n17, B1 => n58, B2 => n16, ZN => 
                           n104);
   U168 : OAI221_X1 port map( B1 => n97, B2 => n18, C1 => n1, C2 => n19, A => 
                           n155, ZN => n120);
   U169 : AOI22_X1 port map( A1 => A(27), A2 => n100, B1 => A(26), B2 => n101, 
                           ZN => n155);
   U170 : AOI221_X1 port map( B1 => n60, B2 => A(13), C1 => n59, C2 => A(12), A
                           => n156, ZN => n108);
   U171 : OAI22_X1 port map( A1 => n43, A2 => n58, B1 => n45, B2 => n57, ZN => 
                           n156);
   U172 : OAI221_X1 port map( B1 => n89, B2 => n92, C1 => n132, C2 => n9, A => 
                           n157, ZN => B(0));
   U173 : AOI222_X1 port map( A1 => n68, A2 => n73, B1 => n55, B2 => n158, C1 
                           => n66, C2 => n44, ZN => n157);
   U174 : AOI221_X1 port map( B1 => n60, B2 => A(11), C1 => n59, C2 => A(10), A
                           => n159, ZN => n70);
   U175 : OAI22_X1 port map( A1 => n46, A2 => n58, B1 => n47, B2 => n57, ZN => 
                           n159);
   U176 : OAI221_X1 port map( B1 => n97, B2 => n52, C1 => n2, C2 => n53, A => 
                           n161, ZN => n158);
   U177 : AOI22_X1 port map( A1 => A(1), A2 => n100, B1 => A(0), B2 => n101, ZN
                           => n161);
   U178 : NAND2_X1 port map( A1 => n56, A2 => n9, ZN => n62);
   U179 : OAI221_X1 port map( B1 => n97, B2 => n37, C1 => n2, C2 => n39, A => 
                           n162, ZN => n73);
   U180 : AOI22_X1 port map( A1 => A(13), A2 => n100, B1 => A(12), B2 => n101, 
                           ZN => n162);
   U181 : AND2_X1 port map( A1 => SH(2), A2 => n160, ZN => n68);
   U182 : NOR2_X1 port map( A1 => n5, A2 => n8, ZN => n160);
   U183 : AOI221_X1 port map( B1 => n75, B2 => n115, C1 => n74, C2 => n56, A =>
                           n10, ZN => n132);
   U184 : AOI22_X1 port map( A1 => n130, A2 => n112, B1 => n118, B2 => n116, ZN
                           => n163);
   U185 : OAI221_X1 port map( B1 => n97, B2 => n20, C1 => n1, C2 => n21, A => 
                           n164, ZN => n116);
   U186 : AOI22_X1 port map( A1 => A(25), A2 => n100, B1 => A(24), B2 => n101, 
                           ZN => n164);
   U187 : NOR2_X1 port map( A1 => n5, A2 => SH(2), ZN => n118);
   U188 : OAI221_X1 port map( B1 => n97, B2 => n16, C1 => n1, C2 => n17, A => 
                           n165, ZN => n112);
   U189 : AOI22_X1 port map( A1 => A(29), A2 => n100, B1 => A(28), B2 => n101, 
                           ZN => n165);
   U190 : NOR2_X1 port map( A1 => n4, A2 => n5, ZN => n130);
   U191 : NAND2_X1 port map( A1 => n4, A2 => n5, ZN => n143);
   U192 : OAI221_X1 port map( B1 => n97, B2 => n30, C1 => n2, C2 => n32, A => 
                           n166, ZN => n74);
   U193 : AOI22_X1 port map( A1 => A(17), A2 => n100, B1 => A(16), B2 => n101, 
                           ZN => n166);
   U194 : OAI221_X1 port map( B1 => n58, B2 => n27, C1 => n29, C2 => n57, A => 
                           n167, ZN => n75);
   U195 : AOI22_X1 port map( A1 => A(23), A2 => n60, B1 => A(22), B2 => n59, ZN
                           => n167);
   U196 : NAND2_X1 port map( A1 => n115, A2 => n9, ZN => n92);
   U197 : NOR2_X1 port map( A1 => n4, A2 => SH(3), ZN => n115);
   U198 : AOI221_X1 port map( B1 => n60, B2 => A(7), C1 => n59, C2 => A(6), A 
                           => n168, ZN => n89);
   U199 : OAI22_X1 port map( A1 => n50, A2 => n58, B1 => n51, B2 => n57, ZN => 
                           n168);
   U200 : NAND2_X1 port map( A1 => SH(1), A2 => n3, ZN => n98);
   U201 : NAND2_X1 port map( A1 => SH(1), A2 => SH(0), ZN => n97);

end SYN_mx2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity SHIFTER_GENERIC_N32_DW_sla_0 is

   port( A : in std_logic_vector (31 downto 0);  SH : in std_logic_vector (4 
         downto 0);  SH_TC : in std_logic;  B : out std_logic_vector (31 downto
         0));

end SHIFTER_GENERIC_N32_DW_sla_0;

architecture SYN_mx2 of SHIFTER_GENERIC_N32_DW_sla_0 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component NOR2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal B_31_port, B_30_port, B_29_port, B_28_port, B_27_port, B_26_port, 
      B_25_port, B_24_port, B_23_port, B_22_port, B_21_port, B_20_port, 
      B_19_port, B_18_port, B_17_port, B_16_port, B_15_port, B_14_port, 
      B_13_port, B_12_port, B_11_port, B_10_port, B_9_port, B_8_port, B_7_port,
      B_6_port, B_5_port, B_4_port, B_3_port, B_2_port, B_1_port, n1, n2, n3, 
      n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19,
      n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34
      , n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, 
      n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63
      , n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, 
      n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92
      , n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, 
      n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116, n117, 
      n118, n119, n120, n121, n122, n123, n124, n125, n126, n127, n128, n129, 
      n130, n131, n132, n133, n134, n135, n136, n137, n138, n139, n140, n141, 
      n142, n143, n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, 
      n154, n155, n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, 
      n166, n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177, 
      n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188 : 
      std_logic;

begin
   B <= ( B_31_port, B_30_port, B_29_port, B_28_port, B_27_port, B_26_port, 
      B_25_port, B_24_port, B_23_port, B_22_port, B_21_port, B_20_port, 
      B_19_port, B_18_port, B_17_port, B_16_port, B_15_port, B_14_port, 
      B_13_port, B_12_port, B_11_port, B_10_port, B_9_port, B_8_port, B_7_port,
      B_6_port, B_5_port, B_4_port, B_3_port, B_2_port, B_1_port, A(0) );
   
   U2 : NOR2_X2 port map( A1 => SH(2), A2 => SH(3), ZN => n130);
   U3 : INV_X1 port map( A => n82, ZN => n72);
   U4 : INV_X1 port map( A => n15, ZN => n18);
   U5 : INV_X1 port map( A => n114, ZN => n73);
   U6 : BUF_X1 port map( A => n94, Z => n10);
   U7 : BUF_X1 port map( A => n94, Z => n11);
   U8 : AND2_X1 port map( A1 => n166, A2 => n14, ZN => n88);
   U9 : BUF_X1 port map( A => n93, Z => n7);
   U10 : BUF_X1 port map( A => n93, Z => n8);
   U11 : BUF_X1 port map( A => n90, Z => n1);
   U12 : BUF_X1 port map( A => n90, Z => n2);
   U13 : BUF_X1 port map( A => n91, Z => n4);
   U14 : BUF_X1 port map( A => n91, Z => n5);
   U15 : BUF_X1 port map( A => SH(4), Z => n15);
   U16 : BUF_X1 port map( A => SH(4), Z => n16);
   U17 : BUF_X1 port map( A => n93, Z => n9);
   U18 : BUF_X1 port map( A => n94, Z => n12);
   U19 : BUF_X1 port map( A => n90, Z => n3);
   U20 : BUF_X1 port map( A => n91, Z => n6);
   U21 : BUF_X1 port map( A => SH(4), Z => n17);
   U22 : INV_X1 port map( A => n168, ZN => n55);
   U23 : INV_X1 port map( A => n171, ZN => n58);
   U24 : INV_X1 port map( A => n177, ZN => n60);
   U25 : INV_X1 port map( A => n181, ZN => n62);
   U26 : INV_X1 port map( A => n185, ZN => n65);
   U27 : INV_X1 port map( A => n131, ZN => n67);
   U28 : INV_X1 port map( A => n173, ZN => n48);
   U29 : INV_X1 port map( A => n75, ZN => n70);
   U30 : INV_X1 port map( A => n153, ZN => n69);
   U31 : INV_X1 port map( A => n86, ZN => n38);
   U32 : INV_X1 port map( A => n97, ZN => n40);
   U33 : INV_X1 port map( A => n104, ZN => n42);
   U34 : INV_X1 port map( A => n110, ZN => n44);
   U35 : INV_X1 port map( A => n138, ZN => n50);
   U36 : INV_X1 port map( A => n89, ZN => n30);
   U37 : INV_X1 port map( A => n99, ZN => n32);
   U38 : INV_X1 port map( A => n106, ZN => n34);
   U39 : INV_X1 port map( A => n112, ZN => n36);
   U40 : NAND2_X1 port map( A1 => n17, A2 => A(0), ZN => n75);
   U41 : INV_X1 port map( A => A(29), ZN => n19);
   U42 : INV_X1 port map( A => n186, ZN => n66);
   U43 : INV_X1 port map( A => A(12), ZN => n49);
   U44 : INV_X1 port map( A => A(23), ZN => n29);
   U45 : INV_X1 port map( A => A(14), ZN => n46);
   U46 : INV_X1 port map( A => A(17), ZN => n41);
   U47 : INV_X1 port map( A => A(21), ZN => n33);
   U48 : INV_X1 port map( A => A(13), ZN => n47);
   U49 : INV_X1 port map( A => A(22), ZN => n31);
   U50 : INV_X1 port map( A => A(16), ZN => n43);
   U51 : INV_X1 port map( A => A(15), ZN => n45);
   U52 : INV_X1 port map( A => A(9), ZN => n53);
   U53 : INV_X1 port map( A => A(7), ZN => n56);
   U54 : INV_X1 port map( A => A(10), ZN => n52);
   U55 : INV_X1 port map( A => A(11), ZN => n51);
   U56 : INV_X1 port map( A => A(8), ZN => n54);
   U57 : INV_X1 port map( A => A(2), ZN => n64);
   U58 : INV_X1 port map( A => A(28), ZN => n20);
   U59 : INV_X1 port map( A => A(27), ZN => n21);
   U60 : INV_X1 port map( A => A(26), ZN => n23);
   U61 : INV_X1 port map( A => A(25), ZN => n25);
   U62 : INV_X1 port map( A => A(24), ZN => n27);
   U63 : INV_X1 port map( A => A(3), ZN => n63);
   U64 : INV_X1 port map( A => A(18), ZN => n39);
   U65 : INV_X1 port map( A => A(0), ZN => n71);
   U66 : INV_X1 port map( A => A(4), ZN => n61);
   U67 : INV_X1 port map( A => A(6), ZN => n57);
   U68 : INV_X1 port map( A => A(19), ZN => n37);
   U69 : INV_X1 port map( A => A(20), ZN => n35);
   U70 : INV_X1 port map( A => A(1), ZN => n68);
   U71 : INV_X1 port map( A => A(5), ZN => n59);
   U72 : INV_X1 port map( A => n118, ZN => n22);
   U73 : INV_X1 port map( A => n123, ZN => n24);
   U74 : INV_X1 port map( A => n135, ZN => n26);
   U75 : INV_X1 port map( A => n141, ZN => n28);
   U76 : INV_X1 port map( A => SH(0), ZN => n13);
   U77 : INV_X1 port map( A => SH(2), ZN => n14);
   U78 : OAI21_X1 port map( B1 => n15, B2 => n74, A => n75, ZN => B_9_port);
   U79 : OAI21_X1 port map( B1 => n15, B2 => n76, A => n75, ZN => B_8_port);
   U80 : OAI21_X1 port map( B1 => n15, B2 => n77, A => n75, ZN => B_7_port);
   U81 : OAI21_X1 port map( B1 => n15, B2 => n78, A => n75, ZN => B_6_port);
   U82 : OAI21_X1 port map( B1 => n15, B2 => n79, A => n75, ZN => B_5_port);
   U83 : OAI21_X1 port map( B1 => n16, B2 => n80, A => n75, ZN => B_4_port);
   U84 : OAI21_X1 port map( B1 => n16, B2 => n81, A => n75, ZN => B_3_port);
   U85 : OAI221_X1 port map( B1 => n22, B2 => n82, C1 => n83, C2 => n18, A => 
                           n84, ZN => B_31_port);
   U86 : AOI222_X1 port map( A1 => n85, A2 => n86, B1 => n73, B2 => n87, C1 => 
                           n88, C2 => n89, ZN => n84);
   U87 : OAI221_X1 port map( B1 => n2, B2 => n19, C1 => n5, C2 => n20, A => n92
                           , ZN => n87);
   U88 : AOI22_X1 port map( A1 => A(30), A2 => n8, B1 => A(31), B2 => n11, ZN 
                           => n92);
   U89 : OAI221_X1 port map( B1 => n24, B2 => n82, C1 => n95, C2 => n18, A => 
                           n96, ZN => B_30_port);
   U90 : AOI222_X1 port map( A1 => n85, A2 => n97, B1 => n73, B2 => n98, C1 => 
                           n88, C2 => n99, ZN => n96);
   U91 : OAI221_X1 port map( B1 => n1, B2 => n20, C1 => n4, C2 => n21, A => 
                           n100, ZN => n98);
   U92 : AOI22_X1 port map( A1 => A(29), A2 => n7, B1 => A(30), B2 => n10, ZN 
                           => n100);
   U93 : OAI21_X1 port map( B1 => n16, B2 => n101, A => n75, ZN => B_2_port);
   U94 : OAI221_X1 port map( B1 => n26, B2 => n82, C1 => n102, C2 => n18, A => 
                           n103, ZN => B_29_port);
   U95 : AOI222_X1 port map( A1 => n85, A2 => n104, B1 => n73, B2 => n105, C1 
                           => n88, C2 => n106, ZN => n103);
   U96 : OAI221_X1 port map( B1 => n1, B2 => n21, C1 => n4, C2 => n23, A => 
                           n107, ZN => n105);
   U97 : AOI22_X1 port map( A1 => A(28), A2 => n7, B1 => A(29), B2 => n10, ZN 
                           => n107);
   U98 : OAI221_X1 port map( B1 => n28, B2 => n82, C1 => n108, C2 => n18, A => 
                           n109, ZN => B_28_port);
   U99 : AOI222_X1 port map( A1 => n85, A2 => n110, B1 => n73, B2 => n111, C1 
                           => n88, C2 => n112, ZN => n109);
   U100 : OAI221_X1 port map( B1 => n1, B2 => n23, C1 => n4, C2 => n25, A => 
                           n113, ZN => n111);
   U101 : AOI22_X1 port map( A1 => A(27), A2 => n7, B1 => A(28), B2 => n10, ZN 
                           => n113);
   U102 : OAI221_X1 port map( B1 => n22, B2 => n114, C1 => n115, C2 => n18, A 
                           => n116, ZN => B_27_port);
   U103 : AOI222_X1 port map( A1 => n72, A2 => n89, B1 => n88, B2 => n86, C1 =>
                           n85, C2 => n117, ZN => n116);
   U104 : OAI221_X1 port map( B1 => n1, B2 => n25, C1 => n4, C2 => n27, A => 
                           n119, ZN => n118);
   U105 : AOI22_X1 port map( A1 => A(26), A2 => n7, B1 => A(27), B2 => n10, ZN 
                           => n119);
   U106 : OAI221_X1 port map( B1 => n24, B2 => n114, C1 => n120, C2 => n18, A 
                           => n121, ZN => B_26_port);
   U107 : AOI222_X1 port map( A1 => n72, A2 => n99, B1 => n88, B2 => n97, C1 =>
                           n85, C2 => n122, ZN => n121);
   U108 : OAI221_X1 port map( B1 => n1, B2 => n27, C1 => n4, C2 => n29, A => 
                           n124, ZN => n123);
   U109 : AOI22_X1 port map( A1 => A(25), A2 => n7, B1 => A(26), B2 => n10, ZN 
                           => n124);
   U110 : OAI221_X1 port map( B1 => n26, B2 => n114, C1 => n74, C2 => n18, A =>
                           n125, ZN => B_25_port);
   U111 : AOI222_X1 port map( A1 => n72, A2 => n106, B1 => n88, B2 => n104, C1 
                           => n85, C2 => n126, ZN => n125);
   U112 : AOI221_X1 port map( B1 => n127, B2 => n128, C1 => n129, C2 => n130, A
                           => n67, ZN => n74);
   U113 : AOI21_X1 port map( B1 => n132, B2 => n133, A => n134, ZN => n131);
   U114 : OAI221_X1 port map( B1 => n1, B2 => n29, C1 => n4, C2 => n31, A => 
                           n136, ZN => n135);
   U115 : AOI22_X1 port map( A1 => A(24), A2 => n7, B1 => A(25), B2 => n10, ZN 
                           => n136);
   U116 : OAI221_X1 port map( B1 => n28, B2 => n114, C1 => n76, C2 => n18, A =>
                           n137, ZN => B_24_port);
   U117 : AOI222_X1 port map( A1 => n72, A2 => n112, B1 => n88, B2 => n110, C1 
                           => n85, C2 => n138, ZN => n137);
   U118 : AOI221_X1 port map( B1 => n139, B2 => n128, C1 => n140, C2 => n130, A
                           => n69, ZN => n76);
   U119 : OAI221_X1 port map( B1 => n1, B2 => n31, C1 => n4, C2 => n33, A => 
                           n142, ZN => n141);
   U120 : AOI22_X1 port map( A1 => A(23), A2 => n7, B1 => A(24), B2 => n10, ZN 
                           => n142);
   U121 : OAI221_X1 port map( B1 => n30, B2 => n114, C1 => n77, C2 => n18, A =>
                           n143, ZN => B_23_port);
   U122 : AOI222_X1 port map( A1 => n72, A2 => n86, B1 => n88, B2 => n117, C1 
                           => n85, C2 => n144, ZN => n143);
   U123 : AOI221_X1 port map( B1 => n145, B2 => n128, C1 => n146, C2 => n130, A
                           => n69, ZN => n77);
   U124 : OAI221_X1 port map( B1 => n1, B2 => n33, C1 => n4, C2 => n35, A => 
                           n147, ZN => n89);
   U125 : AOI22_X1 port map( A1 => A(22), A2 => n7, B1 => A(23), B2 => n10, ZN 
                           => n147);
   U126 : OAI221_X1 port map( B1 => n32, B2 => n114, C1 => n78, C2 => n18, A =>
                           n148, ZN => B_22_port);
   U127 : AOI222_X1 port map( A1 => n72, A2 => n97, B1 => n88, B2 => n122, C1 
                           => n85, C2 => n149, ZN => n148);
   U128 : AOI221_X1 port map( B1 => n66, B2 => n128, C1 => n150, C2 => n130, A 
                           => n69, ZN => n78);
   U129 : OAI221_X1 port map( B1 => n1, B2 => n35, C1 => n5, C2 => n37, A => 
                           n151, ZN => n99);
   U130 : AOI22_X1 port map( A1 => A(21), A2 => n7, B1 => A(22), B2 => n10, ZN 
                           => n151);
   U131 : OAI221_X1 port map( B1 => n34, B2 => n114, C1 => n79, C2 => n18, A =>
                           n152, ZN => B_21_port);
   U132 : AOI222_X1 port map( A1 => n72, A2 => n104, B1 => n88, B2 => n126, C1 
                           => n85, C2 => n129, ZN => n152);
   U133 : AOI221_X1 port map( B1 => n133, B2 => n128, C1 => n127, C2 => n130, A
                           => n69, ZN => n79);
   U134 : OAI221_X1 port map( B1 => n1, B2 => n37, C1 => n5, C2 => n39, A => 
                           n154, ZN => n106);
   U135 : AOI22_X1 port map( A1 => A(20), A2 => n7, B1 => A(21), B2 => n10, ZN 
                           => n154);
   U136 : OAI221_X1 port map( B1 => n36, B2 => n114, C1 => n80, C2 => n18, A =>
                           n155, ZN => B_20_port);
   U137 : AOI222_X1 port map( A1 => n72, A2 => n110, B1 => n88, B2 => n138, C1 
                           => n85, C2 => n140, ZN => n155);
   U138 : AOI21_X1 port map( B1 => n139, B2 => n130, A => n156, ZN => n80);
   U139 : OAI221_X1 port map( B1 => n1, B2 => n39, C1 => n5, C2 => n41, A => 
                           n157, ZN => n112);
   U140 : AOI22_X1 port map( A1 => A(19), A2 => n7, B1 => A(20), B2 => n11, ZN 
                           => n157);
   U141 : OAI21_X1 port map( B1 => n16, B2 => n158, A => n75, ZN => B_1_port);
   U142 : OAI221_X1 port map( B1 => n38, B2 => n114, C1 => n81, C2 => n18, A =>
                           n159, ZN => B_19_port);
   U143 : AOI222_X1 port map( A1 => n72, A2 => n117, B1 => n88, B2 => n144, C1 
                           => n85, C2 => n146, ZN => n159);
   U144 : AOI21_X1 port map( B1 => n145, B2 => n130, A => n156, ZN => n81);
   U145 : OAI221_X1 port map( B1 => n2, B2 => n41, C1 => n5, C2 => n43, A => 
                           n160, ZN => n86);
   U146 : AOI22_X1 port map( A1 => A(18), A2 => n8, B1 => A(19), B2 => n11, ZN 
                           => n160);
   U147 : OAI221_X1 port map( B1 => n40, B2 => n114, C1 => n101, C2 => n18, A 
                           => n161, ZN => B_18_port);
   U148 : AOI222_X1 port map( A1 => n72, A2 => n122, B1 => n88, B2 => n149, C1 
                           => n85, C2 => n150, ZN => n161);
   U149 : AOI21_X1 port map( B1 => n66, B2 => n130, A => n156, ZN => n101);
   U150 : OAI221_X1 port map( B1 => n2, B2 => n43, C1 => n5, C2 => n45, A => 
                           n162, ZN => n97);
   U151 : AOI22_X1 port map( A1 => A(17), A2 => n8, B1 => A(18), B2 => n11, ZN 
                           => n162);
   U152 : OAI221_X1 port map( B1 => n42, B2 => n114, C1 => n158, C2 => n18, A 
                           => n163, ZN => B_17_port);
   U153 : AOI222_X1 port map( A1 => n72, A2 => n126, B1 => n88, B2 => n129, C1 
                           => n85, C2 => n127, ZN => n163);
   U154 : AOI21_X1 port map( B1 => n133, B2 => n130, A => n156, ZN => n158);
   U155 : OAI21_X1 port map( B1 => n71, B2 => n14, A => n153, ZN => n156);
   U156 : OAI221_X1 port map( B1 => n2, B2 => n45, C1 => n5, C2 => n46, A => 
                           n164, ZN => n104);
   U157 : AOI22_X1 port map( A1 => A(16), A2 => n8, B1 => A(17), B2 => n11, ZN 
                           => n164);
   U158 : OAI221_X1 port map( B1 => n50, B2 => n82, C1 => n44, C2 => n114, A =>
                           n165, ZN => B_16_port);
   U159 : AOI221_X1 port map( B1 => n85, B2 => n139, C1 => n88, C2 => n140, A 
                           => n70, ZN => n165);
   U160 : AND2_X1 port map( A1 => n166, A2 => SH(2), ZN => n85);
   U161 : AND2_X1 port map( A1 => SH(3), A2 => n18, ZN => n166);
   U162 : NAND2_X1 port map( A1 => n130, A2 => n18, ZN => n114);
   U163 : OAI221_X1 port map( B1 => n2, B2 => n46, C1 => n5, C2 => n47, A => 
                           n167, ZN => n110);
   U164 : AOI22_X1 port map( A1 => A(15), A2 => n8, B1 => A(16), B2 => n11, ZN 
                           => n167);
   U165 : NAND2_X1 port map( A1 => n128, A2 => n18, ZN => n82);
   U166 : OAI21_X1 port map( B1 => n16, B2 => n83, A => n75, ZN => B_15_port);
   U167 : AOI221_X1 port map( B1 => n144, B2 => n128, C1 => n117, C2 => n130, A
                           => n55, ZN => n83);
   U168 : AOI22_X1 port map( A1 => n169, A2 => n145, B1 => n132, B2 => n146, ZN
                           => n168);
   U169 : OAI221_X1 port map( B1 => n2, B2 => n47, C1 => n5, C2 => n49, A => 
                           n170, ZN => n117);
   U170 : AOI22_X1 port map( A1 => A(14), A2 => n8, B1 => A(15), B2 => n11, ZN 
                           => n170);
   U171 : OAI21_X1 port map( B1 => n16, B2 => n95, A => n75, ZN => B_14_port);
   U172 : AOI221_X1 port map( B1 => n149, B2 => n128, C1 => n122, C2 => n130, A
                           => n58, ZN => n95);
   U173 : AOI22_X1 port map( A1 => n169, A2 => n66, B1 => n132, B2 => n150, ZN 
                           => n171);
   U174 : OAI221_X1 port map( B1 => n2, B2 => n49, C1 => n5, C2 => n51, A => 
                           n172, ZN => n122);
   U175 : AOI22_X1 port map( A1 => A(13), A2 => n8, B1 => A(14), B2 => n11, ZN 
                           => n172);
   U176 : OAI21_X1 port map( B1 => n16, B2 => n102, A => n75, ZN => B_13_port);
   U177 : AOI221_X1 port map( B1 => n133, B2 => n169, C1 => n127, C2 => n132, A
                           => n48, ZN => n102);
   U178 : AOI22_X1 port map( A1 => n128, A2 => n129, B1 => n130, B2 => n126, ZN
                           => n173);
   U179 : OAI221_X1 port map( B1 => n2, B2 => n51, C1 => n5, C2 => n52, A => 
                           n174, ZN => n126);
   U180 : AOI22_X1 port map( A1 => A(12), A2 => n8, B1 => A(13), B2 => n11, ZN 
                           => n174);
   U181 : OAI221_X1 port map( B1 => n2, B2 => n56, C1 => n5, C2 => n57, A => 
                           n175, ZN => n129);
   U182 : AOI22_X1 port map( A1 => A(8), A2 => n8, B1 => A(9), B2 => n11, ZN =>
                           n175);
   U183 : OAI221_X1 port map( B1 => n2, B2 => n63, C1 => n6, C2 => n64, A => 
                           n176, ZN => n127);
   U184 : AOI22_X1 port map( A1 => A(4), A2 => n8, B1 => A(5), B2 => n11, ZN =>
                           n176);
   U185 : AND2_X1 port map( A1 => SH(2), A2 => SH(3), ZN => n169);
   U186 : MUX2_X1 port map( A => A(0), B => A(1), S => n10, Z => n133);
   U187 : OAI21_X1 port map( B1 => n17, B2 => n108, A => n75, ZN => B_12_port);
   U188 : AOI221_X1 port map( B1 => n140, B2 => n128, C1 => n138, C2 => n130, A
                           => n60, ZN => n108);
   U189 : AOI21_X1 port map( B1 => n132, B2 => n139, A => n134, ZN => n177);
   U190 : OAI221_X1 port map( B1 => n2, B2 => n64, C1 => n68, C2 => n4, A => 
                           n178, ZN => n139);
   U191 : AOI22_X1 port map( A1 => n9, A2 => A(3), B1 => A(4), B2 => n11, ZN =>
                           n178);
   U192 : OAI221_X1 port map( B1 => n2, B2 => n52, C1 => n6, C2 => n53, A => 
                           n179, ZN => n138);
   U193 : AOI22_X1 port map( A1 => A(11), A2 => n8, B1 => A(12), B2 => n11, ZN 
                           => n179);
   U194 : OAI221_X1 port map( B1 => n3, B2 => n57, C1 => n6, C2 => n59, A => 
                           n180, ZN => n140);
   U195 : AOI22_X1 port map( A1 => A(7), A2 => n8, B1 => A(8), B2 => n12, ZN =>
                           n180);
   U196 : OAI21_X1 port map( B1 => n17, B2 => n115, A => n75, ZN => B_11_port);
   U197 : AOI221_X1 port map( B1 => n146, B2 => n128, C1 => n144, C2 => n130, A
                           => n62, ZN => n115);
   U198 : AOI21_X1 port map( B1 => n132, B2 => n145, A => n134, ZN => n181);
   U199 : OAI221_X1 port map( B1 => n68, B2 => n3, C1 => n71, C2 => n4, A => 
                           n182, ZN => n145);
   U200 : AOI22_X1 port map( A1 => n9, A2 => A(2), B1 => A(3), B2 => n12, ZN =>
                           n182);
   U201 : OAI221_X1 port map( B1 => n3, B2 => n53, C1 => n6, C2 => n54, A => 
                           n183, ZN => n144);
   U202 : AOI22_X1 port map( A1 => A(10), A2 => n9, B1 => A(11), B2 => n12, ZN 
                           => n183);
   U203 : OAI221_X1 port map( B1 => n3, B2 => n59, C1 => n6, C2 => n61, A => 
                           n184, ZN => n146);
   U204 : AOI22_X1 port map( A1 => A(6), A2 => n9, B1 => A(7), B2 => n12, ZN =>
                           n184);
   U205 : OAI21_X1 port map( B1 => n17, B2 => n120, A => n75, ZN => B_10_port);
   U206 : AOI221_X1 port map( B1 => n150, B2 => n128, C1 => n149, C2 => n130, A
                           => n65, ZN => n120);
   U207 : AOI21_X1 port map( B1 => n132, B2 => n66, A => n134, ZN => n185);
   U208 : NOR2_X1 port map( A1 => n14, A2 => n153, ZN => n134);
   U209 : NAND2_X1 port map( A1 => SH(3), A2 => A(0), ZN => n153);
   U210 : AOI222_X1 port map( A1 => n10, A2 => A(2), B1 => A(1), B2 => n9, C1 
                           => A(0), C2 => SH(1), ZN => n186);
   U211 : AND2_X1 port map( A1 => SH(3), A2 => n14, ZN => n132);
   U212 : OAI221_X1 port map( B1 => n3, B2 => n54, C1 => n4, C2 => n56, A => 
                           n187, ZN => n149);
   U213 : AOI22_X1 port map( A1 => A(9), A2 => n9, B1 => A(10), B2 => n12, ZN 
                           => n187);
   U214 : NOR2_X1 port map( A1 => n14, A2 => SH(3), ZN => n128);
   U215 : OAI221_X1 port map( B1 => n1, B2 => n61, C1 => n63, C2 => n4, A => 
                           n188, ZN => n150);
   U216 : AOI22_X1 port map( A1 => A(5), A2 => n7, B1 => A(6), B2 => n10, ZN =>
                           n188);
   U217 : NOR2_X1 port map( A1 => SH(0), A2 => SH(1), ZN => n94);
   U218 : NOR2_X1 port map( A1 => n13, A2 => SH(1), ZN => n93);
   U219 : NAND2_X1 port map( A1 => SH(0), A2 => SH(1), ZN => n91);
   U220 : NAND2_X1 port map( A1 => SH(1), A2 => n13, ZN => n90);

end SYN_mx2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity SHIFTER_GENERIC_N32_DW01_ash_0 is

   port( A : in std_logic_vector (31 downto 0);  DATA_TC : in std_logic;  SH : 
         in std_logic_vector (4 downto 0);  SH_TC : in std_logic;  B : out 
         std_logic_vector (31 downto 0));

end SHIFTER_GENERIC_N32_DW01_ash_0;

architecture SYN_mx2 of SHIFTER_GENERIC_N32_DW01_ash_0 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   signal ML_int_1_31_port, ML_int_1_30_port, ML_int_1_29_port, 
      ML_int_1_28_port, ML_int_1_27_port, ML_int_1_26_port, ML_int_1_25_port, 
      ML_int_1_24_port, ML_int_1_23_port, ML_int_1_22_port, ML_int_1_21_port, 
      ML_int_1_20_port, ML_int_1_19_port, ML_int_1_18_port, ML_int_1_17_port, 
      ML_int_1_16_port, ML_int_1_15_port, ML_int_1_14_port, ML_int_1_13_port, 
      ML_int_1_12_port, ML_int_1_11_port, ML_int_1_10_port, ML_int_1_9_port, 
      ML_int_1_8_port, ML_int_1_7_port, ML_int_1_6_port, ML_int_1_5_port, 
      ML_int_1_4_port, ML_int_1_3_port, ML_int_1_2_port, ML_int_1_1_port, 
      ML_int_1_0_port, ML_int_2_31_port, ML_int_2_30_port, ML_int_2_29_port, 
      ML_int_2_28_port, ML_int_2_27_port, ML_int_2_26_port, ML_int_2_25_port, 
      ML_int_2_24_port, ML_int_2_23_port, ML_int_2_22_port, ML_int_2_21_port, 
      ML_int_2_20_port, ML_int_2_19_port, ML_int_2_18_port, ML_int_2_17_port, 
      ML_int_2_16_port, ML_int_2_15_port, ML_int_2_14_port, ML_int_2_13_port, 
      ML_int_2_12_port, ML_int_2_11_port, ML_int_2_10_port, ML_int_2_9_port, 
      ML_int_2_8_port, ML_int_2_7_port, ML_int_2_6_port, ML_int_2_5_port, 
      ML_int_2_4_port, ML_int_2_3_port, ML_int_2_2_port, ML_int_2_1_port, 
      ML_int_2_0_port, ML_int_3_31_port, ML_int_3_30_port, ML_int_3_29_port, 
      ML_int_3_28_port, ML_int_3_27_port, ML_int_3_26_port, ML_int_3_25_port, 
      ML_int_3_24_port, ML_int_3_23_port, ML_int_3_22_port, ML_int_3_21_port, 
      ML_int_3_20_port, ML_int_3_19_port, ML_int_3_18_port, ML_int_3_17_port, 
      ML_int_3_16_port, ML_int_3_15_port, ML_int_3_14_port, ML_int_3_13_port, 
      ML_int_3_12_port, ML_int_3_11_port, ML_int_3_10_port, ML_int_3_9_port, 
      ML_int_3_8_port, ML_int_3_7_port, ML_int_3_6_port, ML_int_3_5_port, 
      ML_int_3_4_port, ML_int_3_3_port, ML_int_3_2_port, ML_int_3_1_port, 
      ML_int_3_0_port, ML_int_4_31_port, ML_int_4_30_port, ML_int_4_29_port, 
      ML_int_4_28_port, ML_int_4_27_port, ML_int_4_26_port, ML_int_4_25_port, 
      ML_int_4_24_port, ML_int_4_23_port, ML_int_4_22_port, ML_int_4_21_port, 
      ML_int_4_20_port, ML_int_4_19_port, ML_int_4_18_port, ML_int_4_17_port, 
      ML_int_4_16_port, ML_int_4_15_port, ML_int_4_14_port, ML_int_4_13_port, 
      ML_int_4_12_port, ML_int_4_11_port, ML_int_4_10_port, ML_int_4_9_port, 
      ML_int_4_8_port, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, 
      n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28
      : std_logic;

begin
   
   M1_4_31 : MUX2_X1 port map( A => ML_int_4_31_port, B => ML_int_4_15_port, S 
                           => n11, Z => B(31));
   M1_4_30 : MUX2_X1 port map( A => ML_int_4_30_port, B => ML_int_4_14_port, S 
                           => n11, Z => B(30));
   M1_4_29 : MUX2_X1 port map( A => ML_int_4_29_port, B => ML_int_4_13_port, S 
                           => n11, Z => B(29));
   M1_4_28 : MUX2_X1 port map( A => ML_int_4_28_port, B => ML_int_4_12_port, S 
                           => n11, Z => B(28));
   M1_4_27 : MUX2_X1 port map( A => ML_int_4_27_port, B => ML_int_4_11_port, S 
                           => n11, Z => B(27));
   M1_4_26 : MUX2_X1 port map( A => ML_int_4_26_port, B => ML_int_4_10_port, S 
                           => n11, Z => B(26));
   M1_4_25 : MUX2_X1 port map( A => ML_int_4_25_port, B => ML_int_4_9_port, S 
                           => n11, Z => B(25));
   M1_4_24 : MUX2_X1 port map( A => ML_int_4_24_port, B => ML_int_4_8_port, S 
                           => n11, Z => B(24));
   M1_4_23 : MUX2_X1 port map( A => ML_int_4_23_port, B => n13, S => n11, Z => 
                           B(23));
   M1_4_22 : MUX2_X1 port map( A => ML_int_4_22_port, B => n14, S => n11, Z => 
                           B(22));
   M1_4_21 : MUX2_X1 port map( A => ML_int_4_21_port, B => n15, S => n11, Z => 
                           B(21));
   M1_4_20 : MUX2_X1 port map( A => ML_int_4_20_port, B => n16, S => n11, Z => 
                           B(20));
   M1_4_19 : MUX2_X1 port map( A => ML_int_4_19_port, B => n17, S => SH(4), Z 
                           => B(19));
   M1_4_18 : MUX2_X1 port map( A => ML_int_4_18_port, B => n18, S => n11, Z => 
                           B(18));
   M1_4_17 : MUX2_X1 port map( A => ML_int_4_17_port, B => n19, S => SH(4), Z 
                           => B(17));
   M1_4_16 : MUX2_X1 port map( A => ML_int_4_16_port, B => n20, S => SH(4), Z 
                           => B(16));
   M1_3_31 : MUX2_X1 port map( A => ML_int_3_31_port, B => ML_int_3_23_port, S 
                           => n9, Z => ML_int_4_31_port);
   M1_3_30 : MUX2_X1 port map( A => ML_int_3_30_port, B => ML_int_3_22_port, S 
                           => n9, Z => ML_int_4_30_port);
   M1_3_29 : MUX2_X1 port map( A => ML_int_3_29_port, B => ML_int_3_21_port, S 
                           => n9, Z => ML_int_4_29_port);
   M1_3_28 : MUX2_X1 port map( A => ML_int_3_28_port, B => ML_int_3_20_port, S 
                           => n9, Z => ML_int_4_28_port);
   M1_3_27 : MUX2_X1 port map( A => ML_int_3_27_port, B => ML_int_3_19_port, S 
                           => n9, Z => ML_int_4_27_port);
   M1_3_26 : MUX2_X1 port map( A => ML_int_3_26_port, B => ML_int_3_18_port, S 
                           => n9, Z => ML_int_4_26_port);
   M1_3_25 : MUX2_X1 port map( A => ML_int_3_25_port, B => ML_int_3_17_port, S 
                           => n9, Z => ML_int_4_25_port);
   M1_3_24 : MUX2_X1 port map( A => ML_int_3_24_port, B => ML_int_3_16_port, S 
                           => n9, Z => ML_int_4_24_port);
   M1_3_23 : MUX2_X1 port map( A => ML_int_3_23_port, B => ML_int_3_15_port, S 
                           => n9, Z => ML_int_4_23_port);
   M1_3_22 : MUX2_X1 port map( A => ML_int_3_22_port, B => ML_int_3_14_port, S 
                           => n9, Z => ML_int_4_22_port);
   M1_3_21 : MUX2_X1 port map( A => ML_int_3_21_port, B => ML_int_3_13_port, S 
                           => SH(3), Z => ML_int_4_21_port);
   M1_3_20 : MUX2_X1 port map( A => ML_int_3_20_port, B => ML_int_3_12_port, S 
                           => n9, Z => ML_int_4_20_port);
   M1_3_19 : MUX2_X1 port map( A => ML_int_3_19_port, B => ML_int_3_11_port, S 
                           => n9, Z => ML_int_4_19_port);
   M1_3_18 : MUX2_X1 port map( A => ML_int_3_18_port, B => ML_int_3_10_port, S 
                           => n9, Z => ML_int_4_18_port);
   M1_3_17 : MUX2_X1 port map( A => ML_int_3_17_port, B => ML_int_3_9_port, S 
                           => n9, Z => ML_int_4_17_port);
   M1_3_16 : MUX2_X1 port map( A => ML_int_3_16_port, B => ML_int_3_8_port, S 
                           => n9, Z => ML_int_4_16_port);
   M1_3_15 : MUX2_X1 port map( A => ML_int_3_15_port, B => ML_int_3_7_port, S 
                           => n9, Z => ML_int_4_15_port);
   M1_3_14 : MUX2_X1 port map( A => ML_int_3_14_port, B => ML_int_3_6_port, S 
                           => n9, Z => ML_int_4_14_port);
   M1_3_13 : MUX2_X1 port map( A => ML_int_3_13_port, B => ML_int_3_5_port, S 
                           => n9, Z => ML_int_4_13_port);
   M1_3_12 : MUX2_X1 port map( A => ML_int_3_12_port, B => ML_int_3_4_port, S 
                           => n9, Z => ML_int_4_12_port);
   M1_3_11 : MUX2_X1 port map( A => ML_int_3_11_port, B => ML_int_3_3_port, S 
                           => n9, Z => ML_int_4_11_port);
   M1_3_10 : MUX2_X1 port map( A => ML_int_3_10_port, B => ML_int_3_2_port, S 
                           => n9, Z => ML_int_4_10_port);
   M1_3_9 : MUX2_X1 port map( A => ML_int_3_9_port, B => ML_int_3_1_port, S => 
                           n9, Z => ML_int_4_9_port);
   M1_3_8 : MUX2_X1 port map( A => ML_int_3_8_port, B => ML_int_3_0_port, S => 
                           n9, Z => ML_int_4_8_port);
   M1_2_31 : MUX2_X1 port map( A => ML_int_2_31_port, B => ML_int_2_27_port, S 
                           => n7, Z => ML_int_3_31_port);
   M1_2_30 : MUX2_X1 port map( A => ML_int_2_30_port, B => ML_int_2_26_port, S 
                           => n7, Z => ML_int_3_30_port);
   M1_2_29 : MUX2_X1 port map( A => ML_int_2_29_port, B => ML_int_2_25_port, S 
                           => n7, Z => ML_int_3_29_port);
   M1_2_28 : MUX2_X1 port map( A => ML_int_2_28_port, B => ML_int_2_24_port, S 
                           => n7, Z => ML_int_3_28_port);
   M1_2_27 : MUX2_X1 port map( A => ML_int_2_27_port, B => ML_int_2_23_port, S 
                           => n7, Z => ML_int_3_27_port);
   M1_2_26 : MUX2_X1 port map( A => ML_int_2_26_port, B => ML_int_2_22_port, S 
                           => n7, Z => ML_int_3_26_port);
   M1_2_25 : MUX2_X1 port map( A => ML_int_2_25_port, B => ML_int_2_21_port, S 
                           => SH(2), Z => ML_int_3_25_port);
   M1_2_24 : MUX2_X1 port map( A => ML_int_2_24_port, B => ML_int_2_20_port, S 
                           => n7, Z => ML_int_3_24_port);
   M1_2_23 : MUX2_X1 port map( A => ML_int_2_23_port, B => ML_int_2_19_port, S 
                           => SH(2), Z => ML_int_3_23_port);
   M1_2_22 : MUX2_X1 port map( A => ML_int_2_22_port, B => ML_int_2_18_port, S 
                           => n7, Z => ML_int_3_22_port);
   M1_2_21 : MUX2_X1 port map( A => ML_int_2_21_port, B => ML_int_2_17_port, S 
                           => SH(2), Z => ML_int_3_21_port);
   M1_2_20 : MUX2_X1 port map( A => ML_int_2_20_port, B => ML_int_2_16_port, S 
                           => n7, Z => ML_int_3_20_port);
   M1_2_19 : MUX2_X1 port map( A => ML_int_2_19_port, B => ML_int_2_15_port, S 
                           => SH(2), Z => ML_int_3_19_port);
   M1_2_18 : MUX2_X1 port map( A => ML_int_2_18_port, B => ML_int_2_14_port, S 
                           => n7, Z => ML_int_3_18_port);
   M1_2_17 : MUX2_X1 port map( A => ML_int_2_17_port, B => ML_int_2_13_port, S 
                           => SH(2), Z => ML_int_3_17_port);
   M1_2_16 : MUX2_X1 port map( A => ML_int_2_16_port, B => ML_int_2_12_port, S 
                           => n7, Z => ML_int_3_16_port);
   M1_2_15 : MUX2_X1 port map( A => ML_int_2_15_port, B => ML_int_2_11_port, S 
                           => n7, Z => ML_int_3_15_port);
   M1_2_14 : MUX2_X1 port map( A => ML_int_2_14_port, B => ML_int_2_10_port, S 
                           => n7, Z => ML_int_3_14_port);
   M1_2_13 : MUX2_X1 port map( A => ML_int_2_13_port, B => ML_int_2_9_port, S 
                           => n7, Z => ML_int_3_13_port);
   M1_2_12 : MUX2_X1 port map( A => ML_int_2_12_port, B => ML_int_2_8_port, S 
                           => n7, Z => ML_int_3_12_port);
   M1_2_11 : MUX2_X1 port map( A => ML_int_2_11_port, B => ML_int_2_7_port, S 
                           => n7, Z => ML_int_3_11_port);
   M1_2_10 : MUX2_X1 port map( A => ML_int_2_10_port, B => ML_int_2_6_port, S 
                           => n7, Z => ML_int_3_10_port);
   M1_2_9 : MUX2_X1 port map( A => ML_int_2_9_port, B => ML_int_2_5_port, S => 
                           n7, Z => ML_int_3_9_port);
   M1_2_8 : MUX2_X1 port map( A => ML_int_2_8_port, B => ML_int_2_4_port, S => 
                           n7, Z => ML_int_3_8_port);
   M1_2_7 : MUX2_X1 port map( A => ML_int_2_7_port, B => ML_int_2_3_port, S => 
                           n7, Z => ML_int_3_7_port);
   M1_2_6 : MUX2_X1 port map( A => ML_int_2_6_port, B => ML_int_2_2_port, S => 
                           n7, Z => ML_int_3_6_port);
   M1_2_5 : MUX2_X1 port map( A => ML_int_2_5_port, B => ML_int_2_1_port, S => 
                           n7, Z => ML_int_3_5_port);
   M1_2_4 : MUX2_X1 port map( A => ML_int_2_4_port, B => ML_int_2_0_port, S => 
                           n7, Z => ML_int_3_4_port);
   M1_1_31 : MUX2_X1 port map( A => ML_int_1_31_port, B => ML_int_1_29_port, S 
                           => n5, Z => ML_int_2_31_port);
   M1_1_30 : MUX2_X1 port map( A => ML_int_1_30_port, B => ML_int_1_28_port, S 
                           => n4, Z => ML_int_2_30_port);
   M1_1_29 : MUX2_X1 port map( A => ML_int_1_29_port, B => ML_int_1_27_port, S 
                           => n5, Z => ML_int_2_29_port);
   M1_1_28 : MUX2_X1 port map( A => ML_int_1_28_port, B => ML_int_1_26_port, S 
                           => n4, Z => ML_int_2_28_port);
   M1_1_27 : MUX2_X1 port map( A => ML_int_1_27_port, B => ML_int_1_25_port, S 
                           => n5, Z => ML_int_2_27_port);
   M1_1_26 : MUX2_X1 port map( A => ML_int_1_26_port, B => ML_int_1_24_port, S 
                           => n4, Z => ML_int_2_26_port);
   M1_1_25 : MUX2_X1 port map( A => ML_int_1_25_port, B => ML_int_1_23_port, S 
                           => n5, Z => ML_int_2_25_port);
   M1_1_24 : MUX2_X1 port map( A => ML_int_1_24_port, B => ML_int_1_22_port, S 
                           => n5, Z => ML_int_2_24_port);
   M1_1_23 : MUX2_X1 port map( A => ML_int_1_23_port, B => ML_int_1_21_port, S 
                           => n5, Z => ML_int_2_23_port);
   M1_1_22 : MUX2_X1 port map( A => ML_int_1_22_port, B => ML_int_1_20_port, S 
                           => n5, Z => ML_int_2_22_port);
   M1_1_21 : MUX2_X1 port map( A => ML_int_1_21_port, B => ML_int_1_19_port, S 
                           => n5, Z => ML_int_2_21_port);
   M1_1_20 : MUX2_X1 port map( A => ML_int_1_20_port, B => ML_int_1_18_port, S 
                           => n5, Z => ML_int_2_20_port);
   M1_1_19 : MUX2_X1 port map( A => ML_int_1_19_port, B => ML_int_1_17_port, S 
                           => n5, Z => ML_int_2_19_port);
   M1_1_18 : MUX2_X1 port map( A => ML_int_1_18_port, B => ML_int_1_16_port, S 
                           => n5, Z => ML_int_2_18_port);
   M1_1_17 : MUX2_X1 port map( A => ML_int_1_17_port, B => ML_int_1_15_port, S 
                           => n5, Z => ML_int_2_17_port);
   M1_1_16 : MUX2_X1 port map( A => ML_int_1_16_port, B => ML_int_1_14_port, S 
                           => n5, Z => ML_int_2_16_port);
   M1_1_15 : MUX2_X1 port map( A => ML_int_1_15_port, B => ML_int_1_13_port, S 
                           => n5, Z => ML_int_2_15_port);
   M1_1_14 : MUX2_X1 port map( A => ML_int_1_14_port, B => ML_int_1_12_port, S 
                           => n5, Z => ML_int_2_14_port);
   M1_1_13 : MUX2_X1 port map( A => ML_int_1_13_port, B => ML_int_1_11_port, S 
                           => n4, Z => ML_int_2_13_port);
   M1_1_12 : MUX2_X1 port map( A => ML_int_1_12_port, B => ML_int_1_10_port, S 
                           => n4, Z => ML_int_2_12_port);
   M1_1_11 : MUX2_X1 port map( A => ML_int_1_11_port, B => ML_int_1_9_port, S 
                           => n4, Z => ML_int_2_11_port);
   M1_1_10 : MUX2_X1 port map( A => ML_int_1_10_port, B => ML_int_1_8_port, S 
                           => n4, Z => ML_int_2_10_port);
   M1_1_9 : MUX2_X1 port map( A => ML_int_1_9_port, B => ML_int_1_7_port, S => 
                           n4, Z => ML_int_2_9_port);
   M1_1_8 : MUX2_X1 port map( A => ML_int_1_8_port, B => ML_int_1_6_port, S => 
                           n4, Z => ML_int_2_8_port);
   M1_1_7 : MUX2_X1 port map( A => ML_int_1_7_port, B => ML_int_1_5_port, S => 
                           n4, Z => ML_int_2_7_port);
   M1_1_6 : MUX2_X1 port map( A => ML_int_1_6_port, B => ML_int_1_4_port, S => 
                           n4, Z => ML_int_2_6_port);
   M1_1_5 : MUX2_X1 port map( A => ML_int_1_5_port, B => ML_int_1_3_port, S => 
                           n4, Z => ML_int_2_5_port);
   M1_1_4 : MUX2_X1 port map( A => ML_int_1_4_port, B => ML_int_1_2_port, S => 
                           n4, Z => ML_int_2_4_port);
   M1_1_3 : MUX2_X1 port map( A => ML_int_1_3_port, B => ML_int_1_1_port, S => 
                           n4, Z => ML_int_2_3_port);
   M1_1_2 : MUX2_X1 port map( A => ML_int_1_2_port, B => ML_int_1_0_port, S => 
                           n4, Z => ML_int_2_2_port);
   M1_0_31 : MUX2_X1 port map( A => A(31), B => A(30), S => n2, Z => 
                           ML_int_1_31_port);
   M1_0_30 : MUX2_X1 port map( A => A(30), B => A(29), S => n1, Z => 
                           ML_int_1_30_port);
   M1_0_29 : MUX2_X1 port map( A => A(29), B => A(28), S => n2, Z => 
                           ML_int_1_29_port);
   M1_0_28 : MUX2_X1 port map( A => A(28), B => A(27), S => n1, Z => 
                           ML_int_1_28_port);
   M1_0_27 : MUX2_X1 port map( A => A(27), B => A(26), S => n2, Z => 
                           ML_int_1_27_port);
   M1_0_26 : MUX2_X1 port map( A => A(26), B => A(25), S => n1, Z => 
                           ML_int_1_26_port);
   M1_0_25 : MUX2_X1 port map( A => A(25), B => A(24), S => n2, Z => 
                           ML_int_1_25_port);
   M1_0_24 : MUX2_X1 port map( A => A(24), B => A(23), S => n2, Z => 
                           ML_int_1_24_port);
   M1_0_23 : MUX2_X1 port map( A => A(23), B => A(22), S => n2, Z => 
                           ML_int_1_23_port);
   M1_0_22 : MUX2_X1 port map( A => A(22), B => A(21), S => n2, Z => 
                           ML_int_1_22_port);
   M1_0_21 : MUX2_X1 port map( A => A(21), B => A(20), S => n2, Z => 
                           ML_int_1_21_port);
   M1_0_20 : MUX2_X1 port map( A => A(20), B => A(19), S => n2, Z => 
                           ML_int_1_20_port);
   M1_0_19 : MUX2_X1 port map( A => A(19), B => A(18), S => n2, Z => 
                           ML_int_1_19_port);
   M1_0_18 : MUX2_X1 port map( A => A(18), B => A(17), S => n2, Z => 
                           ML_int_1_18_port);
   M1_0_17 : MUX2_X1 port map( A => A(17), B => A(16), S => n2, Z => 
                           ML_int_1_17_port);
   M1_0_16 : MUX2_X1 port map( A => A(16), B => A(15), S => n2, Z => 
                           ML_int_1_16_port);
   M1_0_15 : MUX2_X1 port map( A => A(15), B => A(14), S => n2, Z => 
                           ML_int_1_15_port);
   M1_0_14 : MUX2_X1 port map( A => A(14), B => A(13), S => n2, Z => 
                           ML_int_1_14_port);
   M1_0_13 : MUX2_X1 port map( A => A(13), B => A(12), S => n2, Z => 
                           ML_int_1_13_port);
   M1_0_12 : MUX2_X1 port map( A => A(12), B => A(11), S => n1, Z => 
                           ML_int_1_12_port);
   M1_0_11 : MUX2_X1 port map( A => A(11), B => A(10), S => n1, Z => 
                           ML_int_1_11_port);
   M1_0_10 : MUX2_X1 port map( A => A(10), B => A(9), S => n1, Z => 
                           ML_int_1_10_port);
   M1_0_9 : MUX2_X1 port map( A => A(9), B => A(8), S => n1, Z => 
                           ML_int_1_9_port);
   M1_0_8 : MUX2_X1 port map( A => A(8), B => A(7), S => n1, Z => 
                           ML_int_1_8_port);
   M1_0_7 : MUX2_X1 port map( A => A(7), B => A(6), S => n1, Z => 
                           ML_int_1_7_port);
   M1_0_6 : MUX2_X1 port map( A => A(6), B => A(5), S => n1, Z => 
                           ML_int_1_6_port);
   M1_0_5 : MUX2_X1 port map( A => A(5), B => A(4), S => n1, Z => 
                           ML_int_1_5_port);
   M1_0_4 : MUX2_X1 port map( A => A(4), B => A(3), S => n1, Z => 
                           ML_int_1_4_port);
   M1_0_3 : MUX2_X1 port map( A => A(3), B => A(2), S => n1, Z => 
                           ML_int_1_3_port);
   M1_0_2 : MUX2_X1 port map( A => A(2), B => A(1), S => n1, Z => 
                           ML_int_1_2_port);
   M1_0_1 : MUX2_X1 port map( A => A(1), B => A(0), S => n1, Z => 
                           ML_int_1_1_port);
   U3 : INV_X1 port map( A => n12, ZN => n11);
   U4 : INV_X1 port map( A => n21, ZN => n13);
   U5 : INV_X1 port map( A => n22, ZN => n14);
   U6 : INV_X1 port map( A => n23, ZN => n15);
   U7 : INV_X1 port map( A => n24, ZN => n16);
   U8 : INV_X1 port map( A => n25, ZN => n17);
   U9 : INV_X1 port map( A => n26, ZN => n18);
   U10 : INV_X1 port map( A => n27, ZN => n19);
   U11 : INV_X1 port map( A => n28, ZN => n20);
   U12 : INV_X1 port map( A => n8, ZN => n7);
   U13 : INV_X1 port map( A => n6, ZN => n5);
   U14 : INV_X1 port map( A => n6, ZN => n4);
   U15 : INV_X1 port map( A => n3, ZN => n2);
   U16 : INV_X1 port map( A => n3, ZN => n1);
   U17 : INV_X1 port map( A => SH(1), ZN => n6);
   U18 : INV_X1 port map( A => SH(0), ZN => n3);
   U19 : INV_X1 port map( A => SH(3), ZN => n10);
   U20 : INV_X1 port map( A => SH(2), ZN => n8);
   U21 : INV_X1 port map( A => n10, ZN => n9);
   U22 : INV_X1 port map( A => SH(4), ZN => n12);
   U23 : AND2_X1 port map( A1 => ML_int_4_9_port, A2 => n12, ZN => B(9));
   U24 : AND2_X1 port map( A1 => ML_int_4_8_port, A2 => n12, ZN => B(8));
   U25 : NOR2_X1 port map( A1 => n11, A2 => n21, ZN => B(7));
   U26 : NOR2_X1 port map( A1 => SH(4), A2 => n22, ZN => B(6));
   U27 : NOR2_X1 port map( A1 => n11, A2 => n23, ZN => B(5));
   U28 : NOR2_X1 port map( A1 => SH(4), A2 => n24, ZN => B(4));
   U29 : NOR2_X1 port map( A1 => n11, A2 => n25, ZN => B(3));
   U30 : NOR2_X1 port map( A1 => SH(4), A2 => n26, ZN => B(2));
   U31 : NOR2_X1 port map( A1 => n11, A2 => n27, ZN => B(1));
   U32 : AND2_X1 port map( A1 => ML_int_4_15_port, A2 => n12, ZN => B(15));
   U33 : AND2_X1 port map( A1 => ML_int_4_14_port, A2 => n12, ZN => B(14));
   U34 : AND2_X1 port map( A1 => ML_int_4_13_port, A2 => n12, ZN => B(13));
   U35 : AND2_X1 port map( A1 => ML_int_4_12_port, A2 => n12, ZN => B(12));
   U36 : AND2_X1 port map( A1 => ML_int_4_11_port, A2 => n12, ZN => B(11));
   U37 : AND2_X1 port map( A1 => ML_int_4_10_port, A2 => n12, ZN => B(10));
   U38 : NOR2_X1 port map( A1 => SH(4), A2 => n28, ZN => B(0));
   U39 : NAND2_X1 port map( A1 => ML_int_3_7_port, A2 => n10, ZN => n21);
   U40 : NAND2_X1 port map( A1 => ML_int_3_6_port, A2 => n10, ZN => n22);
   U41 : NAND2_X1 port map( A1 => ML_int_3_5_port, A2 => n10, ZN => n23);
   U42 : NAND2_X1 port map( A1 => ML_int_3_4_port, A2 => n10, ZN => n24);
   U43 : NAND2_X1 port map( A1 => ML_int_3_3_port, A2 => n10, ZN => n25);
   U44 : NAND2_X1 port map( A1 => ML_int_3_2_port, A2 => n10, ZN => n26);
   U45 : NAND2_X1 port map( A1 => ML_int_3_1_port, A2 => n10, ZN => n27);
   U46 : NAND2_X1 port map( A1 => ML_int_3_0_port, A2 => n10, ZN => n28);
   U47 : AND2_X1 port map( A1 => ML_int_2_3_port, A2 => n8, ZN => 
                           ML_int_3_3_port);
   U48 : AND2_X1 port map( A1 => ML_int_2_2_port, A2 => n8, ZN => 
                           ML_int_3_2_port);
   U49 : AND2_X1 port map( A1 => ML_int_2_1_port, A2 => n8, ZN => 
                           ML_int_3_1_port);
   U50 : AND2_X1 port map( A1 => ML_int_2_0_port, A2 => n8, ZN => 
                           ML_int_3_0_port);
   U51 : AND2_X1 port map( A1 => ML_int_1_1_port, A2 => n6, ZN => 
                           ML_int_2_1_port);
   U52 : AND2_X1 port map( A1 => ML_int_1_0_port, A2 => n6, ZN => 
                           ML_int_2_0_port);
   U53 : AND2_X1 port map( A1 => A(0), A2 => n3, ZN => ML_int_1_0_port);

end SYN_mx2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity DATAPTH_NBIT32_REG_BIT5_DW01_inc_0 is

   port( A : in std_logic_vector (31 downto 0);  SUM : out std_logic_vector (31
         downto 0));

end DATAPTH_NBIT32_REG_BIT5_DW01_inc_0;

architecture SYN_rpl of DATAPTH_NBIT32_REG_BIT5_DW01_inc_0 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component HA_X1
      port( A, B : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal carry_31_port, carry_30_port, carry_29_port, carry_28_port, 
      carry_27_port, carry_26_port, carry_25_port, carry_24_port, carry_23_port
      , carry_22_port, carry_21_port, carry_20_port, carry_19_port, 
      carry_18_port, carry_17_port, carry_16_port, carry_15_port, carry_14_port
      , carry_13_port, carry_12_port, carry_11_port, carry_10_port, 
      carry_9_port, carry_8_port, carry_7_port, carry_6_port, carry_5_port, 
      carry_4_port, carry_3_port, carry_2_port : std_logic;

begin
   
   U1_1_30 : HA_X1 port map( A => A(30), B => carry_30_port, CO => 
                           carry_31_port, S => SUM(30));
   U1_1_29 : HA_X1 port map( A => A(29), B => carry_29_port, CO => 
                           carry_30_port, S => SUM(29));
   U1_1_28 : HA_X1 port map( A => A(28), B => carry_28_port, CO => 
                           carry_29_port, S => SUM(28));
   U1_1_27 : HA_X1 port map( A => A(27), B => carry_27_port, CO => 
                           carry_28_port, S => SUM(27));
   U1_1_26 : HA_X1 port map( A => A(26), B => carry_26_port, CO => 
                           carry_27_port, S => SUM(26));
   U1_1_25 : HA_X1 port map( A => A(25), B => carry_25_port, CO => 
                           carry_26_port, S => SUM(25));
   U1_1_24 : HA_X1 port map( A => A(24), B => carry_24_port, CO => 
                           carry_25_port, S => SUM(24));
   U1_1_23 : HA_X1 port map( A => A(23), B => carry_23_port, CO => 
                           carry_24_port, S => SUM(23));
   U1_1_22 : HA_X1 port map( A => A(22), B => carry_22_port, CO => 
                           carry_23_port, S => SUM(22));
   U1_1_21 : HA_X1 port map( A => A(21), B => carry_21_port, CO => 
                           carry_22_port, S => SUM(21));
   U1_1_20 : HA_X1 port map( A => A(20), B => carry_20_port, CO => 
                           carry_21_port, S => SUM(20));
   U1_1_19 : HA_X1 port map( A => A(19), B => carry_19_port, CO => 
                           carry_20_port, S => SUM(19));
   U1_1_18 : HA_X1 port map( A => A(18), B => carry_18_port, CO => 
                           carry_19_port, S => SUM(18));
   U1_1_17 : HA_X1 port map( A => A(17), B => carry_17_port, CO => 
                           carry_18_port, S => SUM(17));
   U1_1_16 : HA_X1 port map( A => A(16), B => carry_16_port, CO => 
                           carry_17_port, S => SUM(16));
   U1_1_15 : HA_X1 port map( A => A(15), B => carry_15_port, CO => 
                           carry_16_port, S => SUM(15));
   U1_1_14 : HA_X1 port map( A => A(14), B => carry_14_port, CO => 
                           carry_15_port, S => SUM(14));
   U1_1_13 : HA_X1 port map( A => A(13), B => carry_13_port, CO => 
                           carry_14_port, S => SUM(13));
   U1_1_12 : HA_X1 port map( A => A(12), B => carry_12_port, CO => 
                           carry_13_port, S => SUM(12));
   U1_1_11 : HA_X1 port map( A => A(11), B => carry_11_port, CO => 
                           carry_12_port, S => SUM(11));
   U1_1_10 : HA_X1 port map( A => A(10), B => carry_10_port, CO => 
                           carry_11_port, S => SUM(10));
   U1_1_9 : HA_X1 port map( A => A(9), B => carry_9_port, CO => carry_10_port, 
                           S => SUM(9));
   U1_1_8 : HA_X1 port map( A => A(8), B => carry_8_port, CO => carry_9_port, S
                           => SUM(8));
   U1_1_7 : HA_X1 port map( A => A(7), B => carry_7_port, CO => carry_8_port, S
                           => SUM(7));
   U1_1_6 : HA_X1 port map( A => A(6), B => carry_6_port, CO => carry_7_port, S
                           => SUM(6));
   U1_1_5 : HA_X1 port map( A => A(5), B => carry_5_port, CO => carry_6_port, S
                           => SUM(5));
   U1_1_4 : HA_X1 port map( A => A(4), B => carry_4_port, CO => carry_5_port, S
                           => SUM(4));
   U1_1_3 : HA_X1 port map( A => A(3), B => carry_3_port, CO => carry_4_port, S
                           => SUM(3));
   U1_1_2 : HA_X1 port map( A => A(2), B => carry_2_port, CO => carry_3_port, S
                           => SUM(2));
   U1_1_1 : HA_X1 port map( A => A(1), B => A(0), CO => carry_2_port, S => 
                           SUM(1));
   U1 : INV_X1 port map( A => A(0), ZN => SUM(0));
   U2 : XOR2_X1 port map( A => carry_31_port, B => A(31), Z => SUM(31));

end SYN_rpl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_GENERIC_NBIT4_7 is

   port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (3 downto 0));

end MUX21_GENERIC_NBIT4_7;

architecture SYN_struct of MUX21_GENERIC_NBIT4_7 is

   component MUX21_25
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_26
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_27
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_28
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;

begin
   
   gen1_0 : MUX21_28 port map( A => A(0), B => B(0), S => SEL, Y => Y(0));
   gen1_1 : MUX21_27 port map( A => A(1), B => B(1), S => SEL, Y => Y(1));
   gen1_2 : MUX21_26 port map( A => A(2), B => B(2), S => SEL, Y => Y(2));
   gen1_3 : MUX21_25 port map( A => A(3), B => B(3), S => SEL, Y => Y(3));

end SYN_struct;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_GENERIC_NBIT4_6 is

   port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (3 downto 0));

end MUX21_GENERIC_NBIT4_6;

architecture SYN_struct of MUX21_GENERIC_NBIT4_6 is

   component MUX21_21
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_22
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_23
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_24
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;

begin
   
   gen1_0 : MUX21_24 port map( A => A(0), B => B(0), S => SEL, Y => Y(0));
   gen1_1 : MUX21_23 port map( A => A(1), B => B(1), S => SEL, Y => Y(1));
   gen1_2 : MUX21_22 port map( A => A(2), B => B(2), S => SEL, Y => Y(2));
   gen1_3 : MUX21_21 port map( A => A(3), B => B(3), S => SEL, Y => Y(3));

end SYN_struct;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_GENERIC_NBIT4_5 is

   port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (3 downto 0));

end MUX21_GENERIC_NBIT4_5;

architecture SYN_struct of MUX21_GENERIC_NBIT4_5 is

   component MUX21_17
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_18
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_19
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_20
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;

begin
   
   gen1_0 : MUX21_20 port map( A => A(0), B => B(0), S => SEL, Y => Y(0));
   gen1_1 : MUX21_19 port map( A => A(1), B => B(1), S => SEL, Y => Y(1));
   gen1_2 : MUX21_18 port map( A => A(2), B => B(2), S => SEL, Y => Y(2));
   gen1_3 : MUX21_17 port map( A => A(3), B => B(3), S => SEL, Y => Y(3));

end SYN_struct;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_GENERIC_NBIT4_4 is

   port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (3 downto 0));

end MUX21_GENERIC_NBIT4_4;

architecture SYN_struct of MUX21_GENERIC_NBIT4_4 is

   component MUX21_13
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_14
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_15
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_16
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;

begin
   
   gen1_0 : MUX21_16 port map( A => A(0), B => B(0), S => SEL, Y => Y(0));
   gen1_1 : MUX21_15 port map( A => A(1), B => B(1), S => SEL, Y => Y(1));
   gen1_2 : MUX21_14 port map( A => A(2), B => B(2), S => SEL, Y => Y(2));
   gen1_3 : MUX21_13 port map( A => A(3), B => B(3), S => SEL, Y => Y(3));

end SYN_struct;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_GENERIC_NBIT4_3 is

   port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (3 downto 0));

end MUX21_GENERIC_NBIT4_3;

architecture SYN_struct of MUX21_GENERIC_NBIT4_3 is

   component MUX21_9
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_10
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_11
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_12
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;

begin
   
   gen1_0 : MUX21_12 port map( A => A(0), B => B(0), S => SEL, Y => Y(0));
   gen1_1 : MUX21_11 port map( A => A(1), B => B(1), S => SEL, Y => Y(1));
   gen1_2 : MUX21_10 port map( A => A(2), B => B(2), S => SEL, Y => Y(2));
   gen1_3 : MUX21_9 port map( A => A(3), B => B(3), S => SEL, Y => Y(3));

end SYN_struct;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_GENERIC_NBIT4_2 is

   port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (3 downto 0));

end MUX21_GENERIC_NBIT4_2;

architecture SYN_struct of MUX21_GENERIC_NBIT4_2 is

   component MUX21_5
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_6
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_7
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_8
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;

begin
   
   gen1_0 : MUX21_8 port map( A => A(0), B => B(0), S => SEL, Y => Y(0));
   gen1_1 : MUX21_7 port map( A => A(1), B => B(1), S => SEL, Y => Y(1));
   gen1_2 : MUX21_6 port map( A => A(2), B => B(2), S => SEL, Y => Y(2));
   gen1_3 : MUX21_5 port map( A => A(3), B => B(3), S => SEL, Y => Y(3));

end SYN_struct;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_GENERIC_NBIT4_1 is

   port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (3 downto 0));

end MUX21_GENERIC_NBIT4_1;

architecture SYN_struct of MUX21_GENERIC_NBIT4_1 is

   component MUX21_1
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_2
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_3
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_4
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;

begin
   
   gen1_0 : MUX21_4 port map( A => A(0), B => B(0), S => SEL, Y => Y(0));
   gen1_1 : MUX21_3 port map( A => A(1), B => B(1), S => SEL, Y => Y(1));
   gen1_2 : MUX21_2 port map( A => A(2), B => B(2), S => SEL, Y => Y(2));
   gen1_3 : MUX21_1 port map( A => A(3), B => B(3), S => SEL, Y => Y(3));

end SYN_struct;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity RCA_NBIT4_15 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_NBIT4_15;

architecture SYN_BEHAVIORAL of RCA_NBIT4_15 is

   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal add_1_root_add_52_2_carry_1_port, add_1_root_add_52_2_carry_2_port, 
      add_1_root_add_52_2_carry_3_port : std_logic;

begin
   
   add_1_root_add_52_2_U1_0 : FA_X1 port map( A => A(0), B => B(0), CI => Ci, 
                           CO => add_1_root_add_52_2_carry_1_port, S => S(0));
   add_1_root_add_52_2_U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => 
                           add_1_root_add_52_2_carry_1_port, CO => 
                           add_1_root_add_52_2_carry_2_port, S => S(1));
   add_1_root_add_52_2_U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => 
                           add_1_root_add_52_2_carry_2_port, CO => 
                           add_1_root_add_52_2_carry_3_port, S => S(2));
   add_1_root_add_52_2_U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => 
                           add_1_root_add_52_2_carry_3_port, CO => Co, S => 
                           S(3));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity RCA_NBIT4_14 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_NBIT4_14;

architecture SYN_BEHAVIORAL of RCA_NBIT4_14 is

   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal add_1_root_add_52_2_carry_1_port, add_1_root_add_52_2_carry_2_port, 
      add_1_root_add_52_2_carry_3_port : std_logic;

begin
   
   add_1_root_add_52_2_U1_0 : FA_X1 port map( A => A(0), B => B(0), CI => Ci, 
                           CO => add_1_root_add_52_2_carry_1_port, S => S(0));
   add_1_root_add_52_2_U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => 
                           add_1_root_add_52_2_carry_1_port, CO => 
                           add_1_root_add_52_2_carry_2_port, S => S(1));
   add_1_root_add_52_2_U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => 
                           add_1_root_add_52_2_carry_2_port, CO => 
                           add_1_root_add_52_2_carry_3_port, S => S(2));
   add_1_root_add_52_2_U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => 
                           add_1_root_add_52_2_carry_3_port, CO => Co, S => 
                           S(3));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity RCA_NBIT4_13 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_NBIT4_13;

architecture SYN_BEHAVIORAL of RCA_NBIT4_13 is

   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal add_1_root_add_52_2_carry_1_port, add_1_root_add_52_2_carry_2_port, 
      add_1_root_add_52_2_carry_3_port : std_logic;

begin
   
   add_1_root_add_52_2_U1_0 : FA_X1 port map( A => A(0), B => B(0), CI => Ci, 
                           CO => add_1_root_add_52_2_carry_1_port, S => S(0));
   add_1_root_add_52_2_U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => 
                           add_1_root_add_52_2_carry_1_port, CO => 
                           add_1_root_add_52_2_carry_2_port, S => S(1));
   add_1_root_add_52_2_U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => 
                           add_1_root_add_52_2_carry_2_port, CO => 
                           add_1_root_add_52_2_carry_3_port, S => S(2));
   add_1_root_add_52_2_U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => 
                           add_1_root_add_52_2_carry_3_port, CO => Co, S => 
                           S(3));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity RCA_NBIT4_12 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_NBIT4_12;

architecture SYN_BEHAVIORAL of RCA_NBIT4_12 is

   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal add_1_root_add_52_2_carry_1_port, add_1_root_add_52_2_carry_2_port, 
      add_1_root_add_52_2_carry_3_port : std_logic;

begin
   
   add_1_root_add_52_2_U1_0 : FA_X1 port map( A => A(0), B => B(0), CI => Ci, 
                           CO => add_1_root_add_52_2_carry_1_port, S => S(0));
   add_1_root_add_52_2_U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => 
                           add_1_root_add_52_2_carry_1_port, CO => 
                           add_1_root_add_52_2_carry_2_port, S => S(1));
   add_1_root_add_52_2_U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => 
                           add_1_root_add_52_2_carry_2_port, CO => 
                           add_1_root_add_52_2_carry_3_port, S => S(2));
   add_1_root_add_52_2_U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => 
                           add_1_root_add_52_2_carry_3_port, CO => Co, S => 
                           S(3));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity RCA_NBIT4_11 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_NBIT4_11;

architecture SYN_BEHAVIORAL of RCA_NBIT4_11 is

   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal add_1_root_add_52_2_carry_1_port, add_1_root_add_52_2_carry_2_port, 
      add_1_root_add_52_2_carry_3_port : std_logic;

begin
   
   add_1_root_add_52_2_U1_0 : FA_X1 port map( A => A(0), B => B(0), CI => Ci, 
                           CO => add_1_root_add_52_2_carry_1_port, S => S(0));
   add_1_root_add_52_2_U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => 
                           add_1_root_add_52_2_carry_1_port, CO => 
                           add_1_root_add_52_2_carry_2_port, S => S(1));
   add_1_root_add_52_2_U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => 
                           add_1_root_add_52_2_carry_2_port, CO => 
                           add_1_root_add_52_2_carry_3_port, S => S(2));
   add_1_root_add_52_2_U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => 
                           add_1_root_add_52_2_carry_3_port, CO => Co, S => 
                           S(3));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity RCA_NBIT4_10 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_NBIT4_10;

architecture SYN_BEHAVIORAL of RCA_NBIT4_10 is

   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal add_1_root_add_52_2_carry_1_port, add_1_root_add_52_2_carry_2_port, 
      add_1_root_add_52_2_carry_3_port : std_logic;

begin
   
   add_1_root_add_52_2_U1_0 : FA_X1 port map( A => A(0), B => B(0), CI => Ci, 
                           CO => add_1_root_add_52_2_carry_1_port, S => S(0));
   add_1_root_add_52_2_U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => 
                           add_1_root_add_52_2_carry_1_port, CO => 
                           add_1_root_add_52_2_carry_2_port, S => S(1));
   add_1_root_add_52_2_U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => 
                           add_1_root_add_52_2_carry_2_port, CO => 
                           add_1_root_add_52_2_carry_3_port, S => S(2));
   add_1_root_add_52_2_U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => 
                           add_1_root_add_52_2_carry_3_port, CO => Co, S => 
                           S(3));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity RCA_NBIT4_9 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_NBIT4_9;

architecture SYN_BEHAVIORAL of RCA_NBIT4_9 is

   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal add_1_root_add_52_2_carry_1_port, add_1_root_add_52_2_carry_2_port, 
      add_1_root_add_52_2_carry_3_port : std_logic;

begin
   
   add_1_root_add_52_2_U1_0 : FA_X1 port map( A => A(0), B => B(0), CI => Ci, 
                           CO => add_1_root_add_52_2_carry_1_port, S => S(0));
   add_1_root_add_52_2_U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => 
                           add_1_root_add_52_2_carry_1_port, CO => 
                           add_1_root_add_52_2_carry_2_port, S => S(1));
   add_1_root_add_52_2_U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => 
                           add_1_root_add_52_2_carry_2_port, CO => 
                           add_1_root_add_52_2_carry_3_port, S => S(2));
   add_1_root_add_52_2_U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => 
                           add_1_root_add_52_2_carry_3_port, CO => Co, S => 
                           S(3));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity RCA_NBIT4_8 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_NBIT4_8;

architecture SYN_BEHAVIORAL of RCA_NBIT4_8 is

   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal add_1_root_add_52_2_carry_1_port, add_1_root_add_52_2_carry_2_port, 
      add_1_root_add_52_2_carry_3_port : std_logic;

begin
   
   add_1_root_add_52_2_U1_0 : FA_X1 port map( A => A(0), B => B(0), CI => Ci, 
                           CO => add_1_root_add_52_2_carry_1_port, S => S(0));
   add_1_root_add_52_2_U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => 
                           add_1_root_add_52_2_carry_1_port, CO => 
                           add_1_root_add_52_2_carry_2_port, S => S(1));
   add_1_root_add_52_2_U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => 
                           add_1_root_add_52_2_carry_2_port, CO => 
                           add_1_root_add_52_2_carry_3_port, S => S(2));
   add_1_root_add_52_2_U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => 
                           add_1_root_add_52_2_carry_3_port, CO => Co, S => 
                           S(3));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity RCA_NBIT4_7 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_NBIT4_7;

architecture SYN_BEHAVIORAL of RCA_NBIT4_7 is

   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal add_1_root_add_52_2_carry_1_port, add_1_root_add_52_2_carry_2_port, 
      add_1_root_add_52_2_carry_3_port : std_logic;

begin
   
   add_1_root_add_52_2_U1_0 : FA_X1 port map( A => A(0), B => B(0), CI => Ci, 
                           CO => add_1_root_add_52_2_carry_1_port, S => S(0));
   add_1_root_add_52_2_U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => 
                           add_1_root_add_52_2_carry_1_port, CO => 
                           add_1_root_add_52_2_carry_2_port, S => S(1));
   add_1_root_add_52_2_U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => 
                           add_1_root_add_52_2_carry_2_port, CO => 
                           add_1_root_add_52_2_carry_3_port, S => S(2));
   add_1_root_add_52_2_U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => 
                           add_1_root_add_52_2_carry_3_port, CO => Co, S => 
                           S(3));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity RCA_NBIT4_6 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_NBIT4_6;

architecture SYN_BEHAVIORAL of RCA_NBIT4_6 is

   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal add_1_root_add_52_2_carry_1_port, add_1_root_add_52_2_carry_2_port, 
      add_1_root_add_52_2_carry_3_port : std_logic;

begin
   
   add_1_root_add_52_2_U1_0 : FA_X1 port map( A => A(0), B => B(0), CI => Ci, 
                           CO => add_1_root_add_52_2_carry_1_port, S => S(0));
   add_1_root_add_52_2_U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => 
                           add_1_root_add_52_2_carry_1_port, CO => 
                           add_1_root_add_52_2_carry_2_port, S => S(1));
   add_1_root_add_52_2_U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => 
                           add_1_root_add_52_2_carry_2_port, CO => 
                           add_1_root_add_52_2_carry_3_port, S => S(2));
   add_1_root_add_52_2_U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => 
                           add_1_root_add_52_2_carry_3_port, CO => Co, S => 
                           S(3));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity RCA_NBIT4_5 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_NBIT4_5;

architecture SYN_BEHAVIORAL of RCA_NBIT4_5 is

   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal add_1_root_add_52_2_carry_1_port, add_1_root_add_52_2_carry_2_port, 
      add_1_root_add_52_2_carry_3_port : std_logic;

begin
   
   add_1_root_add_52_2_U1_0 : FA_X1 port map( A => A(0), B => B(0), CI => Ci, 
                           CO => add_1_root_add_52_2_carry_1_port, S => S(0));
   add_1_root_add_52_2_U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => 
                           add_1_root_add_52_2_carry_1_port, CO => 
                           add_1_root_add_52_2_carry_2_port, S => S(1));
   add_1_root_add_52_2_U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => 
                           add_1_root_add_52_2_carry_2_port, CO => 
                           add_1_root_add_52_2_carry_3_port, S => S(2));
   add_1_root_add_52_2_U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => 
                           add_1_root_add_52_2_carry_3_port, CO => Co, S => 
                           S(3));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity RCA_NBIT4_4 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_NBIT4_4;

architecture SYN_BEHAVIORAL of RCA_NBIT4_4 is

   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal add_1_root_add_52_2_carry_1_port, add_1_root_add_52_2_carry_2_port, 
      add_1_root_add_52_2_carry_3_port : std_logic;

begin
   
   add_1_root_add_52_2_U1_0 : FA_X1 port map( A => A(0), B => B(0), CI => Ci, 
                           CO => add_1_root_add_52_2_carry_1_port, S => S(0));
   add_1_root_add_52_2_U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => 
                           add_1_root_add_52_2_carry_1_port, CO => 
                           add_1_root_add_52_2_carry_2_port, S => S(1));
   add_1_root_add_52_2_U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => 
                           add_1_root_add_52_2_carry_2_port, CO => 
                           add_1_root_add_52_2_carry_3_port, S => S(2));
   add_1_root_add_52_2_U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => 
                           add_1_root_add_52_2_carry_3_port, CO => Co, S => 
                           S(3));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity RCA_NBIT4_3 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_NBIT4_3;

architecture SYN_BEHAVIORAL of RCA_NBIT4_3 is

   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal add_1_root_add_52_2_carry_1_port, add_1_root_add_52_2_carry_2_port, 
      add_1_root_add_52_2_carry_3_port : std_logic;

begin
   
   add_1_root_add_52_2_U1_0 : FA_X1 port map( A => A(0), B => B(0), CI => Ci, 
                           CO => add_1_root_add_52_2_carry_1_port, S => S(0));
   add_1_root_add_52_2_U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => 
                           add_1_root_add_52_2_carry_1_port, CO => 
                           add_1_root_add_52_2_carry_2_port, S => S(1));
   add_1_root_add_52_2_U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => 
                           add_1_root_add_52_2_carry_2_port, CO => 
                           add_1_root_add_52_2_carry_3_port, S => S(2));
   add_1_root_add_52_2_U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => 
                           add_1_root_add_52_2_carry_3_port, CO => Co, S => 
                           S(3));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity RCA_NBIT4_2 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_NBIT4_2;

architecture SYN_BEHAVIORAL of RCA_NBIT4_2 is

   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal add_1_root_add_52_2_carry_1_port, add_1_root_add_52_2_carry_2_port, 
      add_1_root_add_52_2_carry_3_port : std_logic;

begin
   
   add_1_root_add_52_2_U1_0 : FA_X1 port map( A => A(0), B => B(0), CI => Ci, 
                           CO => add_1_root_add_52_2_carry_1_port, S => S(0));
   add_1_root_add_52_2_U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => 
                           add_1_root_add_52_2_carry_1_port, CO => 
                           add_1_root_add_52_2_carry_2_port, S => S(1));
   add_1_root_add_52_2_U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => 
                           add_1_root_add_52_2_carry_2_port, CO => 
                           add_1_root_add_52_2_carry_3_port, S => S(2));
   add_1_root_add_52_2_U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => 
                           add_1_root_add_52_2_carry_3_port, CO => Co, S => 
                           S(3));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity RCA_NBIT4_1 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_NBIT4_1;

architecture SYN_BEHAVIORAL of RCA_NBIT4_1 is

   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal add_1_root_add_52_2_carry_1_port, add_1_root_add_52_2_carry_2_port, 
      add_1_root_add_52_2_carry_3_port : std_logic;

begin
   
   add_1_root_add_52_2_U1_0 : FA_X1 port map( A => A(0), B => B(0), CI => Ci, 
                           CO => add_1_root_add_52_2_carry_1_port, S => S(0));
   add_1_root_add_52_2_U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => 
                           add_1_root_add_52_2_carry_1_port, CO => 
                           add_1_root_add_52_2_carry_2_port, S => S(1));
   add_1_root_add_52_2_U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => 
                           add_1_root_add_52_2_carry_2_port, CO => 
                           add_1_root_add_52_2_carry_3_port, S => S(2));
   add_1_root_add_52_2_U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => 
                           add_1_root_add_52_2_carry_3_port, CO => Co, S => 
                           S(3));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity P_42 is

   port( p1, P2 : in std_logic;  Co : out std_logic);

end P_42;

architecture SYN_behave of P_42 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => p1, A2 => P2, ZN => Co);

end SYN_behave;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity P_41 is

   port( p1, P2 : in std_logic;  Co : out std_logic);

end P_41;

architecture SYN_behave of P_41 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => p1, A2 => P2, ZN => Co);

end SYN_behave;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity P_40 is

   port( p1, P2 : in std_logic;  Co : out std_logic);

end P_40;

architecture SYN_behave of P_40 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => p1, A2 => P2, ZN => Co);

end SYN_behave;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity P_39 is

   port( p1, P2 : in std_logic;  Co : out std_logic);

end P_39;

architecture SYN_behave of P_39 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => p1, A2 => P2, ZN => Co);

end SYN_behave;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity P_38 is

   port( p1, P2 : in std_logic;  Co : out std_logic);

end P_38;

architecture SYN_behave of P_38 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => p1, A2 => P2, ZN => Co);

end SYN_behave;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity P_37 is

   port( p1, P2 : in std_logic;  Co : out std_logic);

end P_37;

architecture SYN_behave of P_37 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => p1, A2 => P2, ZN => Co);

end SYN_behave;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity P_36 is

   port( p1, P2 : in std_logic;  Co : out std_logic);

end P_36;

architecture SYN_behave of P_36 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => p1, A2 => P2, ZN => Co);

end SYN_behave;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity P_35 is

   port( p1, P2 : in std_logic;  Co : out std_logic);

end P_35;

architecture SYN_behave of P_35 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => p1, A2 => P2, ZN => Co);

end SYN_behave;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity P_34 is

   port( p1, P2 : in std_logic;  Co : out std_logic);

end P_34;

architecture SYN_behave of P_34 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => p1, A2 => P2, ZN => Co);

end SYN_behave;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity P_33 is

   port( p1, P2 : in std_logic;  Co : out std_logic);

end P_33;

architecture SYN_behave of P_33 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => p1, A2 => P2, ZN => Co);

end SYN_behave;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity P_32 is

   port( p1, P2 : in std_logic;  Co : out std_logic);

end P_32;

architecture SYN_behave of P_32 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => p1, A2 => P2, ZN => Co);

end SYN_behave;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity P_31 is

   port( p1, P2 : in std_logic;  Co : out std_logic);

end P_31;

architecture SYN_behave of P_31 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => p1, A2 => P2, ZN => Co);

end SYN_behave;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity P_30 is

   port( p1, P2 : in std_logic;  Co : out std_logic);

end P_30;

architecture SYN_behave of P_30 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => p1, A2 => P2, ZN => Co);

end SYN_behave;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity P_29 is

   port( p1, P2 : in std_logic;  Co : out std_logic);

end P_29;

architecture SYN_behave of P_29 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => p1, A2 => P2, ZN => Co);

end SYN_behave;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity P_28 is

   port( p1, P2 : in std_logic;  Co : out std_logic);

end P_28;

architecture SYN_behave of P_28 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => p1, A2 => P2, ZN => Co);

end SYN_behave;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity P_27 is

   port( p1, P2 : in std_logic;  Co : out std_logic);

end P_27;

architecture SYN_behave of P_27 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => p1, A2 => P2, ZN => Co);

end SYN_behave;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity P_26 is

   port( p1, P2 : in std_logic;  Co : out std_logic);

end P_26;

architecture SYN_behave of P_26 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => p1, A2 => P2, ZN => Co);

end SYN_behave;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity P_25 is

   port( p1, P2 : in std_logic;  Co : out std_logic);

end P_25;

architecture SYN_behave of P_25 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => p1, A2 => P2, ZN => Co);

end SYN_behave;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity P_24 is

   port( p1, P2 : in std_logic;  Co : out std_logic);

end P_24;

architecture SYN_behave of P_24 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => p1, A2 => P2, ZN => Co);

end SYN_behave;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity P_23 is

   port( p1, P2 : in std_logic;  Co : out std_logic);

end P_23;

architecture SYN_behave of P_23 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => p1, A2 => P2, ZN => Co);

end SYN_behave;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity P_22 is

   port( p1, P2 : in std_logic;  Co : out std_logic);

end P_22;

architecture SYN_behave of P_22 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => p1, A2 => P2, ZN => Co);

end SYN_behave;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity P_21 is

   port( p1, P2 : in std_logic;  Co : out std_logic);

end P_21;

architecture SYN_behave of P_21 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => p1, A2 => P2, ZN => Co);

end SYN_behave;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity P_20 is

   port( p1, P2 : in std_logic;  Co : out std_logic);

end P_20;

architecture SYN_behave of P_20 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => p1, A2 => P2, ZN => Co);

end SYN_behave;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity P_19 is

   port( p1, P2 : in std_logic;  Co : out std_logic);

end P_19;

architecture SYN_behave of P_19 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => p1, A2 => P2, ZN => Co);

end SYN_behave;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity P_18 is

   port( p1, P2 : in std_logic;  Co : out std_logic);

end P_18;

architecture SYN_behave of P_18 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => p1, A2 => P2, ZN => Co);

end SYN_behave;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity P_17 is

   port( p1, P2 : in std_logic;  Co : out std_logic);

end P_17;

architecture SYN_behave of P_17 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => p1, A2 => P2, ZN => Co);

end SYN_behave;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity P_16 is

   port( p1, P2 : in std_logic;  Co : out std_logic);

end P_16;

architecture SYN_behave of P_16 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => p1, A2 => P2, ZN => Co);

end SYN_behave;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity P_15 is

   port( p1, P2 : in std_logic;  Co : out std_logic);

end P_15;

architecture SYN_behave of P_15 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => p1, A2 => P2, ZN => Co);

end SYN_behave;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity P_14 is

   port( p1, P2 : in std_logic;  Co : out std_logic);

end P_14;

architecture SYN_behave of P_14 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => p1, A2 => P2, ZN => Co);

end SYN_behave;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity P_13 is

   port( p1, P2 : in std_logic;  Co : out std_logic);

end P_13;

architecture SYN_behave of P_13 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => p1, A2 => P2, ZN => Co);

end SYN_behave;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity P_12 is

   port( p1, P2 : in std_logic;  Co : out std_logic);

end P_12;

architecture SYN_behave of P_12 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => p1, A2 => P2, ZN => Co);

end SYN_behave;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity P_11 is

   port( p1, P2 : in std_logic;  Co : out std_logic);

end P_11;

architecture SYN_behave of P_11 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => p1, A2 => P2, ZN => Co);

end SYN_behave;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity P_10 is

   port( p1, P2 : in std_logic;  Co : out std_logic);

end P_10;

architecture SYN_behave of P_10 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => p1, A2 => P2, ZN => Co);

end SYN_behave;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity P_9 is

   port( p1, P2 : in std_logic;  Co : out std_logic);

end P_9;

architecture SYN_behave of P_9 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => p1, A2 => P2, ZN => Co);

end SYN_behave;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity P_8 is

   port( p1, P2 : in std_logic;  Co : out std_logic);

end P_8;

architecture SYN_behave of P_8 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => p1, A2 => P2, ZN => Co);

end SYN_behave;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity P_7 is

   port( p1, P2 : in std_logic;  Co : out std_logic);

end P_7;

architecture SYN_behave of P_7 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => p1, A2 => P2, ZN => Co);

end SYN_behave;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity P_6 is

   port( p1, P2 : in std_logic;  Co : out std_logic);

end P_6;

architecture SYN_behave of P_6 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => p1, A2 => P2, ZN => Co);

end SYN_behave;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity P_5 is

   port( p1, P2 : in std_logic;  Co : out std_logic);

end P_5;

architecture SYN_behave of P_5 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => p1, A2 => P2, ZN => Co);

end SYN_behave;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity P_4 is

   port( p1, P2 : in std_logic;  Co : out std_logic);

end P_4;

architecture SYN_behave of P_4 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => p1, A2 => P2, ZN => Co);

end SYN_behave;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity P_3 is

   port( p1, P2 : in std_logic;  Co : out std_logic);

end P_3;

architecture SYN_behave of P_3 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => p1, A2 => P2, ZN => Co);

end SYN_behave;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity P_2 is

   port( p1, P2 : in std_logic;  Co : out std_logic);

end P_2;

architecture SYN_behave of P_2 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => p1, A2 => P2, ZN => Co);

end SYN_behave;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity P_1 is

   port( p1, P2 : in std_logic;  Co : out std_logic);

end P_1;

architecture SYN_behave of P_1 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => p1, A2 => P2, ZN => Co);

end SYN_behave;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity CSB_NBIT4_7 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0));

end CSB_NBIT4_7;

architecture SYN_STRUCTURAL of CSB_NBIT4_7 is

   component MUX21_GENERIC_NBIT4_7
      port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component RCA_NBIT4_13
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCA_NBIT4_14
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, out_rca0_3_port, out_rca0_2_port, 
      out_rca0_1_port, out_rca0_0_port, out_rca1_3_port, out_rca1_2_port, 
      out_rca1_1_port, out_rca1_0_port, n_1020, n_1021 : std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA0 : RCA_NBIT4_14 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), A(0)
                           => A(0), B(3) => B(3), B(2) => B(2), B(1) => B(1), 
                           B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           out_rca0_3_port, S(2) => out_rca0_2_port, S(1) => 
                           out_rca0_1_port, S(0) => out_rca0_0_port, Co => 
                           n_1020);
   RCA1 : RCA_NBIT4_13 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), A(0)
                           => A(0), B(3) => B(3), B(2) => B(2), B(1) => B(1), 
                           B(0) => B(0), Ci => X_Logic1_port, S(3) => 
                           out_rca1_3_port, S(2) => out_rca1_2_port, S(1) => 
                           out_rca1_1_port, S(0) => out_rca1_0_port, Co => 
                           n_1021);
   MUXCin : MUX21_GENERIC_NBIT4_7 port map( A(3) => out_rca1_3_port, A(2) => 
                           out_rca1_2_port, A(1) => out_rca1_1_port, A(0) => 
                           out_rca1_0_port, B(3) => out_rca0_3_port, B(2) => 
                           out_rca0_2_port, B(1) => out_rca0_1_port, B(0) => 
                           out_rca0_0_port, SEL => Ci, Y(3) => S(3), Y(2) => 
                           S(2), Y(1) => S(1), Y(0) => S(0));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity CSB_NBIT4_6 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0));

end CSB_NBIT4_6;

architecture SYN_STRUCTURAL of CSB_NBIT4_6 is

   component MUX21_GENERIC_NBIT4_6
      port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component RCA_NBIT4_11
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCA_NBIT4_12
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, out_rca0_3_port, out_rca0_2_port, 
      out_rca0_1_port, out_rca0_0_port, out_rca1_3_port, out_rca1_2_port, 
      out_rca1_1_port, out_rca1_0_port, n_1022, n_1023 : std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA0 : RCA_NBIT4_12 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), A(0)
                           => A(0), B(3) => B(3), B(2) => B(2), B(1) => B(1), 
                           B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           out_rca0_3_port, S(2) => out_rca0_2_port, S(1) => 
                           out_rca0_1_port, S(0) => out_rca0_0_port, Co => 
                           n_1022);
   RCA1 : RCA_NBIT4_11 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), A(0)
                           => A(0), B(3) => B(3), B(2) => B(2), B(1) => B(1), 
                           B(0) => B(0), Ci => X_Logic1_port, S(3) => 
                           out_rca1_3_port, S(2) => out_rca1_2_port, S(1) => 
                           out_rca1_1_port, S(0) => out_rca1_0_port, Co => 
                           n_1023);
   MUXCin : MUX21_GENERIC_NBIT4_6 port map( A(3) => out_rca1_3_port, A(2) => 
                           out_rca1_2_port, A(1) => out_rca1_1_port, A(0) => 
                           out_rca1_0_port, B(3) => out_rca0_3_port, B(2) => 
                           out_rca0_2_port, B(1) => out_rca0_1_port, B(0) => 
                           out_rca0_0_port, SEL => Ci, Y(3) => S(3), Y(2) => 
                           S(2), Y(1) => S(1), Y(0) => S(0));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity CSB_NBIT4_5 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0));

end CSB_NBIT4_5;

architecture SYN_STRUCTURAL of CSB_NBIT4_5 is

   component MUX21_GENERIC_NBIT4_5
      port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component RCA_NBIT4_9
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCA_NBIT4_10
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, out_rca0_3_port, out_rca0_2_port, 
      out_rca0_1_port, out_rca0_0_port, out_rca1_3_port, out_rca1_2_port, 
      out_rca1_1_port, out_rca1_0_port, n_1024, n_1025 : std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA0 : RCA_NBIT4_10 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), A(0)
                           => A(0), B(3) => B(3), B(2) => B(2), B(1) => B(1), 
                           B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           out_rca0_3_port, S(2) => out_rca0_2_port, S(1) => 
                           out_rca0_1_port, S(0) => out_rca0_0_port, Co => 
                           n_1024);
   RCA1 : RCA_NBIT4_9 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), A(0) 
                           => A(0), B(3) => B(3), B(2) => B(2), B(1) => B(1), 
                           B(0) => B(0), Ci => X_Logic1_port, S(3) => 
                           out_rca1_3_port, S(2) => out_rca1_2_port, S(1) => 
                           out_rca1_1_port, S(0) => out_rca1_0_port, Co => 
                           n_1025);
   MUXCin : MUX21_GENERIC_NBIT4_5 port map( A(3) => out_rca1_3_port, A(2) => 
                           out_rca1_2_port, A(1) => out_rca1_1_port, A(0) => 
                           out_rca1_0_port, B(3) => out_rca0_3_port, B(2) => 
                           out_rca0_2_port, B(1) => out_rca0_1_port, B(0) => 
                           out_rca0_0_port, SEL => Ci, Y(3) => S(3), Y(2) => 
                           S(2), Y(1) => S(1), Y(0) => S(0));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity CSB_NBIT4_4 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0));

end CSB_NBIT4_4;

architecture SYN_STRUCTURAL of CSB_NBIT4_4 is

   component MUX21_GENERIC_NBIT4_4
      port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component RCA_NBIT4_7
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCA_NBIT4_8
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, out_rca0_3_port, out_rca0_2_port, 
      out_rca0_1_port, out_rca0_0_port, out_rca1_3_port, out_rca1_2_port, 
      out_rca1_1_port, out_rca1_0_port, n_1026, n_1027 : std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA0 : RCA_NBIT4_8 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), A(0) 
                           => A(0), B(3) => B(3), B(2) => B(2), B(1) => B(1), 
                           B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           out_rca0_3_port, S(2) => out_rca0_2_port, S(1) => 
                           out_rca0_1_port, S(0) => out_rca0_0_port, Co => 
                           n_1026);
   RCA1 : RCA_NBIT4_7 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), A(0) 
                           => A(0), B(3) => B(3), B(2) => B(2), B(1) => B(1), 
                           B(0) => B(0), Ci => X_Logic1_port, S(3) => 
                           out_rca1_3_port, S(2) => out_rca1_2_port, S(1) => 
                           out_rca1_1_port, S(0) => out_rca1_0_port, Co => 
                           n_1027);
   MUXCin : MUX21_GENERIC_NBIT4_4 port map( A(3) => out_rca1_3_port, A(2) => 
                           out_rca1_2_port, A(1) => out_rca1_1_port, A(0) => 
                           out_rca1_0_port, B(3) => out_rca0_3_port, B(2) => 
                           out_rca0_2_port, B(1) => out_rca0_1_port, B(0) => 
                           out_rca0_0_port, SEL => Ci, Y(3) => S(3), Y(2) => 
                           S(2), Y(1) => S(1), Y(0) => S(0));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity CSB_NBIT4_3 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0));

end CSB_NBIT4_3;

architecture SYN_STRUCTURAL of CSB_NBIT4_3 is

   component MUX21_GENERIC_NBIT4_3
      port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component RCA_NBIT4_5
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCA_NBIT4_6
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, out_rca0_3_port, out_rca0_2_port, 
      out_rca0_1_port, out_rca0_0_port, out_rca1_3_port, out_rca1_2_port, 
      out_rca1_1_port, out_rca1_0_port, n_1028, n_1029 : std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA0 : RCA_NBIT4_6 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), A(0) 
                           => A(0), B(3) => B(3), B(2) => B(2), B(1) => B(1), 
                           B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           out_rca0_3_port, S(2) => out_rca0_2_port, S(1) => 
                           out_rca0_1_port, S(0) => out_rca0_0_port, Co => 
                           n_1028);
   RCA1 : RCA_NBIT4_5 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), A(0) 
                           => A(0), B(3) => B(3), B(2) => B(2), B(1) => B(1), 
                           B(0) => B(0), Ci => X_Logic1_port, S(3) => 
                           out_rca1_3_port, S(2) => out_rca1_2_port, S(1) => 
                           out_rca1_1_port, S(0) => out_rca1_0_port, Co => 
                           n_1029);
   MUXCin : MUX21_GENERIC_NBIT4_3 port map( A(3) => out_rca1_3_port, A(2) => 
                           out_rca1_2_port, A(1) => out_rca1_1_port, A(0) => 
                           out_rca1_0_port, B(3) => out_rca0_3_port, B(2) => 
                           out_rca0_2_port, B(1) => out_rca0_1_port, B(0) => 
                           out_rca0_0_port, SEL => Ci, Y(3) => S(3), Y(2) => 
                           S(2), Y(1) => S(1), Y(0) => S(0));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity CSB_NBIT4_2 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0));

end CSB_NBIT4_2;

architecture SYN_STRUCTURAL of CSB_NBIT4_2 is

   component MUX21_GENERIC_NBIT4_2
      port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component RCA_NBIT4_3
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCA_NBIT4_4
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, out_rca0_3_port, out_rca0_2_port, 
      out_rca0_1_port, out_rca0_0_port, out_rca1_3_port, out_rca1_2_port, 
      out_rca1_1_port, out_rca1_0_port, n_1030, n_1031 : std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA0 : RCA_NBIT4_4 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), A(0) 
                           => A(0), B(3) => B(3), B(2) => B(2), B(1) => B(1), 
                           B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           out_rca0_3_port, S(2) => out_rca0_2_port, S(1) => 
                           out_rca0_1_port, S(0) => out_rca0_0_port, Co => 
                           n_1030);
   RCA1 : RCA_NBIT4_3 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), A(0) 
                           => A(0), B(3) => B(3), B(2) => B(2), B(1) => B(1), 
                           B(0) => B(0), Ci => X_Logic1_port, S(3) => 
                           out_rca1_3_port, S(2) => out_rca1_2_port, S(1) => 
                           out_rca1_1_port, S(0) => out_rca1_0_port, Co => 
                           n_1031);
   MUXCin : MUX21_GENERIC_NBIT4_2 port map( A(3) => out_rca1_3_port, A(2) => 
                           out_rca1_2_port, A(1) => out_rca1_1_port, A(0) => 
                           out_rca1_0_port, B(3) => out_rca0_3_port, B(2) => 
                           out_rca0_2_port, B(1) => out_rca0_1_port, B(0) => 
                           out_rca0_0_port, SEL => Ci, Y(3) => S(3), Y(2) => 
                           S(2), Y(1) => S(1), Y(0) => S(0));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity CSB_NBIT4_1 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0));

end CSB_NBIT4_1;

architecture SYN_STRUCTURAL of CSB_NBIT4_1 is

   component MUX21_GENERIC_NBIT4_1
      port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component RCA_NBIT4_1
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCA_NBIT4_2
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, out_rca0_3_port, out_rca0_2_port, 
      out_rca0_1_port, out_rca0_0_port, out_rca1_3_port, out_rca1_2_port, 
      out_rca1_1_port, out_rca1_0_port, n_1032, n_1033 : std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA0 : RCA_NBIT4_2 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), A(0) 
                           => A(0), B(3) => B(3), B(2) => B(2), B(1) => B(1), 
                           B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           out_rca0_3_port, S(2) => out_rca0_2_port, S(1) => 
                           out_rca0_1_port, S(0) => out_rca0_0_port, Co => 
                           n_1032);
   RCA1 : RCA_NBIT4_1 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), A(0) 
                           => A(0), B(3) => B(3), B(2) => B(2), B(1) => B(1), 
                           B(0) => B(0), Ci => X_Logic1_port, S(3) => 
                           out_rca1_3_port, S(2) => out_rca1_2_port, S(1) => 
                           out_rca1_1_port, S(0) => out_rca1_0_port, Co => 
                           n_1033);
   MUXCin : MUX21_GENERIC_NBIT4_1 port map( A(3) => out_rca1_3_port, A(2) => 
                           out_rca1_2_port, A(1) => out_rca1_1_port, A(0) => 
                           out_rca1_0_port, B(3) => out_rca0_3_port, B(2) => 
                           out_rca0_2_port, B(1) => out_rca0_1_port, B(0) => 
                           out_rca0_0_port, SEL => Ci, Y(3) => S(3), Y(2) => 
                           S(2), Y(1) => S(1), Y(0) => S(0));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity PG_42 is

   port( G1, P1, G2, P2 : in std_logic;  gout, pout : out std_logic);

end PG_42;

architecture SYN_arch of PG_42 is

   component P_42
      port( p1, P2 : in std_logic;  Co : out std_logic);
   end component;
   
   component G_42
      port( G1, P, G2 : in std_logic;  Co : out std_logic);
   end component;

begin
   
   g_comp : G_42 port map( G1 => G1, P => P1, G2 => G2, Co => gout);
   p_comp : P_42 port map( p1 => P1, P2 => P2, Co => pout);

end SYN_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity PG_41 is

   port( G1, P1, G2, P2 : in std_logic;  gout, pout : out std_logic);

end PG_41;

architecture SYN_arch of PG_41 is

   component P_41
      port( p1, P2 : in std_logic;  Co : out std_logic);
   end component;
   
   component G_41
      port( G1, P, G2 : in std_logic;  Co : out std_logic);
   end component;

begin
   
   g_comp : G_41 port map( G1 => G1, P => P1, G2 => G2, Co => gout);
   p_comp : P_41 port map( p1 => P1, P2 => P2, Co => pout);

end SYN_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity PG_40 is

   port( G1, P1, G2, P2 : in std_logic;  gout, pout : out std_logic);

end PG_40;

architecture SYN_arch of PG_40 is

   component P_40
      port( p1, P2 : in std_logic;  Co : out std_logic);
   end component;
   
   component G_40
      port( G1, P, G2 : in std_logic;  Co : out std_logic);
   end component;

begin
   
   g_comp : G_40 port map( G1 => G1, P => P1, G2 => G2, Co => gout);
   p_comp : P_40 port map( p1 => P1, P2 => P2, Co => pout);

end SYN_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity PG_39 is

   port( G1, P1, G2, P2 : in std_logic;  gout, pout : out std_logic);

end PG_39;

architecture SYN_arch of PG_39 is

   component P_39
      port( p1, P2 : in std_logic;  Co : out std_logic);
   end component;
   
   component G_39
      port( G1, P, G2 : in std_logic;  Co : out std_logic);
   end component;

begin
   
   g_comp : G_39 port map( G1 => G1, P => P1, G2 => G2, Co => gout);
   p_comp : P_39 port map( p1 => P1, P2 => P2, Co => pout);

end SYN_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity PG_38 is

   port( G1, P1, G2, P2 : in std_logic;  gout, pout : out std_logic);

end PG_38;

architecture SYN_arch of PG_38 is

   component P_38
      port( p1, P2 : in std_logic;  Co : out std_logic);
   end component;
   
   component G_38
      port( G1, P, G2 : in std_logic;  Co : out std_logic);
   end component;

begin
   
   g_comp : G_38 port map( G1 => G1, P => P1, G2 => G2, Co => gout);
   p_comp : P_38 port map( p1 => P1, P2 => P2, Co => pout);

end SYN_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity PG_37 is

   port( G1, P1, G2, P2 : in std_logic;  gout, pout : out std_logic);

end PG_37;

architecture SYN_arch of PG_37 is

   component P_37
      port( p1, P2 : in std_logic;  Co : out std_logic);
   end component;
   
   component G_37
      port( G1, P, G2 : in std_logic;  Co : out std_logic);
   end component;

begin
   
   g_comp : G_37 port map( G1 => G1, P => P1, G2 => G2, Co => gout);
   p_comp : P_37 port map( p1 => P1, P2 => P2, Co => pout);

end SYN_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity PG_36 is

   port( G1, P1, G2, P2 : in std_logic;  gout, pout : out std_logic);

end PG_36;

architecture SYN_arch of PG_36 is

   component P_36
      port( p1, P2 : in std_logic;  Co : out std_logic);
   end component;
   
   component G_36
      port( G1, P, G2 : in std_logic;  Co : out std_logic);
   end component;

begin
   
   g_comp : G_36 port map( G1 => G1, P => P1, G2 => G2, Co => gout);
   p_comp : P_36 port map( p1 => P1, P2 => P2, Co => pout);

end SYN_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity PG_35 is

   port( G1, P1, G2, P2 : in std_logic;  gout, pout : out std_logic);

end PG_35;

architecture SYN_arch of PG_35 is

   component P_35
      port( p1, P2 : in std_logic;  Co : out std_logic);
   end component;
   
   component G_35
      port( G1, P, G2 : in std_logic;  Co : out std_logic);
   end component;

begin
   
   g_comp : G_35 port map( G1 => G1, P => P1, G2 => G2, Co => gout);
   p_comp : P_35 port map( p1 => P1, P2 => P2, Co => pout);

end SYN_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity PG_34 is

   port( G1, P1, G2, P2 : in std_logic;  gout, pout : out std_logic);

end PG_34;

architecture SYN_arch of PG_34 is

   component P_34
      port( p1, P2 : in std_logic;  Co : out std_logic);
   end component;
   
   component G_34
      port( G1, P, G2 : in std_logic;  Co : out std_logic);
   end component;

begin
   
   g_comp : G_34 port map( G1 => G1, P => P1, G2 => G2, Co => gout);
   p_comp : P_34 port map( p1 => P1, P2 => P2, Co => pout);

end SYN_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity PG_33 is

   port( G1, P1, G2, P2 : in std_logic;  gout, pout : out std_logic);

end PG_33;

architecture SYN_arch of PG_33 is

   component P_33
      port( p1, P2 : in std_logic;  Co : out std_logic);
   end component;
   
   component G_33
      port( G1, P, G2 : in std_logic;  Co : out std_logic);
   end component;

begin
   
   g_comp : G_33 port map( G1 => G1, P => P1, G2 => G2, Co => gout);
   p_comp : P_33 port map( p1 => P1, P2 => P2, Co => pout);

end SYN_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity PG_32 is

   port( G1, P1, G2, P2 : in std_logic;  gout, pout : out std_logic);

end PG_32;

architecture SYN_arch of PG_32 is

   component P_32
      port( p1, P2 : in std_logic;  Co : out std_logic);
   end component;
   
   component G_32
      port( G1, P, G2 : in std_logic;  Co : out std_logic);
   end component;

begin
   
   g_comp : G_32 port map( G1 => G1, P => P1, G2 => G2, Co => gout);
   p_comp : P_32 port map( p1 => P1, P2 => P2, Co => pout);

end SYN_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity PG_31 is

   port( G1, P1, G2, P2 : in std_logic;  gout, pout : out std_logic);

end PG_31;

architecture SYN_arch of PG_31 is

   component P_31
      port( p1, P2 : in std_logic;  Co : out std_logic);
   end component;
   
   component G_31
      port( G1, P, G2 : in std_logic;  Co : out std_logic);
   end component;

begin
   
   g_comp : G_31 port map( G1 => G1, P => P1, G2 => G2, Co => gout);
   p_comp : P_31 port map( p1 => P1, P2 => P2, Co => pout);

end SYN_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity PG_30 is

   port( G1, P1, G2, P2 : in std_logic;  gout, pout : out std_logic);

end PG_30;

architecture SYN_arch of PG_30 is

   component P_30
      port( p1, P2 : in std_logic;  Co : out std_logic);
   end component;
   
   component G_30
      port( G1, P, G2 : in std_logic;  Co : out std_logic);
   end component;

begin
   
   g_comp : G_30 port map( G1 => G1, P => P1, G2 => G2, Co => gout);
   p_comp : P_30 port map( p1 => P1, P2 => P2, Co => pout);

end SYN_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity PG_29 is

   port( G1, P1, G2, P2 : in std_logic;  gout, pout : out std_logic);

end PG_29;

architecture SYN_arch of PG_29 is

   component P_29
      port( p1, P2 : in std_logic;  Co : out std_logic);
   end component;
   
   component G_29
      port( G1, P, G2 : in std_logic;  Co : out std_logic);
   end component;

begin
   
   g_comp : G_29 port map( G1 => G1, P => P1, G2 => G2, Co => gout);
   p_comp : P_29 port map( p1 => P1, P2 => P2, Co => pout);

end SYN_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity PG_28 is

   port( G1, P1, G2, P2 : in std_logic;  gout, pout : out std_logic);

end PG_28;

architecture SYN_arch of PG_28 is

   component P_28
      port( p1, P2 : in std_logic;  Co : out std_logic);
   end component;
   
   component G_28
      port( G1, P, G2 : in std_logic;  Co : out std_logic);
   end component;

begin
   
   g_comp : G_28 port map( G1 => G1, P => P1, G2 => G2, Co => gout);
   p_comp : P_28 port map( p1 => P1, P2 => P2, Co => pout);

end SYN_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity PG_27 is

   port( G1, P1, G2, P2 : in std_logic;  gout, pout : out std_logic);

end PG_27;

architecture SYN_arch of PG_27 is

   component P_27
      port( p1, P2 : in std_logic;  Co : out std_logic);
   end component;
   
   component G_27
      port( G1, P, G2 : in std_logic;  Co : out std_logic);
   end component;

begin
   
   g_comp : G_27 port map( G1 => G1, P => P1, G2 => G2, Co => gout);
   p_comp : P_27 port map( p1 => P1, P2 => P2, Co => pout);

end SYN_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity PG_26 is

   port( G1, P1, G2, P2 : in std_logic;  gout, pout : out std_logic);

end PG_26;

architecture SYN_arch of PG_26 is

   component P_26
      port( p1, P2 : in std_logic;  Co : out std_logic);
   end component;
   
   component G_26
      port( G1, P, G2 : in std_logic;  Co : out std_logic);
   end component;

begin
   
   g_comp : G_26 port map( G1 => G1, P => P1, G2 => G2, Co => gout);
   p_comp : P_26 port map( p1 => P1, P2 => P2, Co => pout);

end SYN_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity PG_25 is

   port( G1, P1, G2, P2 : in std_logic;  gout, pout : out std_logic);

end PG_25;

architecture SYN_arch of PG_25 is

   component P_25
      port( p1, P2 : in std_logic;  Co : out std_logic);
   end component;
   
   component G_25
      port( G1, P, G2 : in std_logic;  Co : out std_logic);
   end component;

begin
   
   g_comp : G_25 port map( G1 => G1, P => P1, G2 => G2, Co => gout);
   p_comp : P_25 port map( p1 => P1, P2 => P2, Co => pout);

end SYN_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity PG_24 is

   port( G1, P1, G2, P2 : in std_logic;  gout, pout : out std_logic);

end PG_24;

architecture SYN_arch of PG_24 is

   component P_24
      port( p1, P2 : in std_logic;  Co : out std_logic);
   end component;
   
   component G_24
      port( G1, P, G2 : in std_logic;  Co : out std_logic);
   end component;

begin
   
   g_comp : G_24 port map( G1 => G1, P => P1, G2 => G2, Co => gout);
   p_comp : P_24 port map( p1 => P1, P2 => P2, Co => pout);

end SYN_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity PG_23 is

   port( G1, P1, G2, P2 : in std_logic;  gout, pout : out std_logic);

end PG_23;

architecture SYN_arch of PG_23 is

   component P_23
      port( p1, P2 : in std_logic;  Co : out std_logic);
   end component;
   
   component G_23
      port( G1, P, G2 : in std_logic;  Co : out std_logic);
   end component;

begin
   
   g_comp : G_23 port map( G1 => G1, P => P1, G2 => G2, Co => gout);
   p_comp : P_23 port map( p1 => P1, P2 => P2, Co => pout);

end SYN_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity PG_22 is

   port( G1, P1, G2, P2 : in std_logic;  gout, pout : out std_logic);

end PG_22;

architecture SYN_arch of PG_22 is

   component P_22
      port( p1, P2 : in std_logic;  Co : out std_logic);
   end component;
   
   component G_22
      port( G1, P, G2 : in std_logic;  Co : out std_logic);
   end component;

begin
   
   g_comp : G_22 port map( G1 => G1, P => P1, G2 => G2, Co => gout);
   p_comp : P_22 port map( p1 => P1, P2 => P2, Co => pout);

end SYN_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity PG_21 is

   port( G1, P1, G2, P2 : in std_logic;  gout, pout : out std_logic);

end PG_21;

architecture SYN_arch of PG_21 is

   component P_21
      port( p1, P2 : in std_logic;  Co : out std_logic);
   end component;
   
   component G_21
      port( G1, P, G2 : in std_logic;  Co : out std_logic);
   end component;

begin
   
   g_comp : G_21 port map( G1 => G1, P => P1, G2 => G2, Co => gout);
   p_comp : P_21 port map( p1 => P1, P2 => P2, Co => pout);

end SYN_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity PG_20 is

   port( G1, P1, G2, P2 : in std_logic;  gout, pout : out std_logic);

end PG_20;

architecture SYN_arch of PG_20 is

   component P_20
      port( p1, P2 : in std_logic;  Co : out std_logic);
   end component;
   
   component G_20
      port( G1, P, G2 : in std_logic;  Co : out std_logic);
   end component;

begin
   
   g_comp : G_20 port map( G1 => G1, P => P1, G2 => G2, Co => gout);
   p_comp : P_20 port map( p1 => P1, P2 => P2, Co => pout);

end SYN_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity PG_19 is

   port( G1, P1, G2, P2 : in std_logic;  gout, pout : out std_logic);

end PG_19;

architecture SYN_arch of PG_19 is

   component P_19
      port( p1, P2 : in std_logic;  Co : out std_logic);
   end component;
   
   component G_19
      port( G1, P, G2 : in std_logic;  Co : out std_logic);
   end component;

begin
   
   g_comp : G_19 port map( G1 => G1, P => P1, G2 => G2, Co => gout);
   p_comp : P_19 port map( p1 => P1, P2 => P2, Co => pout);

end SYN_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity PG_18 is

   port( G1, P1, G2, P2 : in std_logic;  gout, pout : out std_logic);

end PG_18;

architecture SYN_arch of PG_18 is

   component P_18
      port( p1, P2 : in std_logic;  Co : out std_logic);
   end component;
   
   component G_18
      port( G1, P, G2 : in std_logic;  Co : out std_logic);
   end component;

begin
   
   g_comp : G_18 port map( G1 => G1, P => P1, G2 => G2, Co => gout);
   p_comp : P_18 port map( p1 => P1, P2 => P2, Co => pout);

end SYN_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity PG_17 is

   port( G1, P1, G2, P2 : in std_logic;  gout, pout : out std_logic);

end PG_17;

architecture SYN_arch of PG_17 is

   component P_17
      port( p1, P2 : in std_logic;  Co : out std_logic);
   end component;
   
   component G_17
      port( G1, P, G2 : in std_logic;  Co : out std_logic);
   end component;

begin
   
   g_comp : G_17 port map( G1 => G1, P => P1, G2 => G2, Co => gout);
   p_comp : P_17 port map( p1 => P1, P2 => P2, Co => pout);

end SYN_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity PG_16 is

   port( G1, P1, G2, P2 : in std_logic;  gout, pout : out std_logic);

end PG_16;

architecture SYN_arch of PG_16 is

   component P_16
      port( p1, P2 : in std_logic;  Co : out std_logic);
   end component;
   
   component G_16
      port( G1, P, G2 : in std_logic;  Co : out std_logic);
   end component;

begin
   
   g_comp : G_16 port map( G1 => G1, P => P1, G2 => G2, Co => gout);
   p_comp : P_16 port map( p1 => P1, P2 => P2, Co => pout);

end SYN_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity PG_15 is

   port( G1, P1, G2, P2 : in std_logic;  gout, pout : out std_logic);

end PG_15;

architecture SYN_arch of PG_15 is

   component P_15
      port( p1, P2 : in std_logic;  Co : out std_logic);
   end component;
   
   component G_15
      port( G1, P, G2 : in std_logic;  Co : out std_logic);
   end component;

begin
   
   g_comp : G_15 port map( G1 => G1, P => P1, G2 => G2, Co => gout);
   p_comp : P_15 port map( p1 => P1, P2 => P2, Co => pout);

end SYN_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity PG_14 is

   port( G1, P1, G2, P2 : in std_logic;  gout, pout : out std_logic);

end PG_14;

architecture SYN_arch of PG_14 is

   component P_14
      port( p1, P2 : in std_logic;  Co : out std_logic);
   end component;
   
   component G_14
      port( G1, P, G2 : in std_logic;  Co : out std_logic);
   end component;

begin
   
   g_comp : G_14 port map( G1 => G1, P => P1, G2 => G2, Co => gout);
   p_comp : P_14 port map( p1 => P1, P2 => P2, Co => pout);

end SYN_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity PG_13 is

   port( G1, P1, G2, P2 : in std_logic;  gout, pout : out std_logic);

end PG_13;

architecture SYN_arch of PG_13 is

   component P_13
      port( p1, P2 : in std_logic;  Co : out std_logic);
   end component;
   
   component G_13
      port( G1, P, G2 : in std_logic;  Co : out std_logic);
   end component;

begin
   
   g_comp : G_13 port map( G1 => G1, P => P1, G2 => G2, Co => gout);
   p_comp : P_13 port map( p1 => P1, P2 => P2, Co => pout);

end SYN_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity PG_12 is

   port( G1, P1, G2, P2 : in std_logic;  gout, pout : out std_logic);

end PG_12;

architecture SYN_arch of PG_12 is

   component P_12
      port( p1, P2 : in std_logic;  Co : out std_logic);
   end component;
   
   component G_12
      port( G1, P, G2 : in std_logic;  Co : out std_logic);
   end component;

begin
   
   g_comp : G_12 port map( G1 => G1, P => P1, G2 => G2, Co => gout);
   p_comp : P_12 port map( p1 => P1, P2 => P2, Co => pout);

end SYN_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity PG_11 is

   port( G1, P1, G2, P2 : in std_logic;  gout, pout : out std_logic);

end PG_11;

architecture SYN_arch of PG_11 is

   component P_11
      port( p1, P2 : in std_logic;  Co : out std_logic);
   end component;
   
   component G_11
      port( G1, P, G2 : in std_logic;  Co : out std_logic);
   end component;

begin
   
   g_comp : G_11 port map( G1 => G1, P => P1, G2 => G2, Co => gout);
   p_comp : P_11 port map( p1 => P1, P2 => P2, Co => pout);

end SYN_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity PG_10 is

   port( G1, P1, G2, P2 : in std_logic;  gout, pout : out std_logic);

end PG_10;

architecture SYN_arch of PG_10 is

   component P_10
      port( p1, P2 : in std_logic;  Co : out std_logic);
   end component;
   
   component G_10
      port( G1, P, G2 : in std_logic;  Co : out std_logic);
   end component;

begin
   
   g_comp : G_10 port map( G1 => G1, P => P1, G2 => G2, Co => gout);
   p_comp : P_10 port map( p1 => P1, P2 => P2, Co => pout);

end SYN_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity PG_9 is

   port( G1, P1, G2, P2 : in std_logic;  gout, pout : out std_logic);

end PG_9;

architecture SYN_arch of PG_9 is

   component P_9
      port( p1, P2 : in std_logic;  Co : out std_logic);
   end component;
   
   component G_9
      port( G1, P, G2 : in std_logic;  Co : out std_logic);
   end component;

begin
   
   g_comp : G_9 port map( G1 => G1, P => P1, G2 => G2, Co => gout);
   p_comp : P_9 port map( p1 => P1, P2 => P2, Co => pout);

end SYN_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity PG_8 is

   port( G1, P1, G2, P2 : in std_logic;  gout, pout : out std_logic);

end PG_8;

architecture SYN_arch of PG_8 is

   component P_8
      port( p1, P2 : in std_logic;  Co : out std_logic);
   end component;
   
   component G_8
      port( G1, P, G2 : in std_logic;  Co : out std_logic);
   end component;

begin
   
   g_comp : G_8 port map( G1 => G1, P => P1, G2 => G2, Co => gout);
   p_comp : P_8 port map( p1 => P1, P2 => P2, Co => pout);

end SYN_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity PG_7 is

   port( G1, P1, G2, P2 : in std_logic;  gout, pout : out std_logic);

end PG_7;

architecture SYN_arch of PG_7 is

   component P_7
      port( p1, P2 : in std_logic;  Co : out std_logic);
   end component;
   
   component G_7
      port( G1, P, G2 : in std_logic;  Co : out std_logic);
   end component;

begin
   
   g_comp : G_7 port map( G1 => G1, P => P1, G2 => G2, Co => gout);
   p_comp : P_7 port map( p1 => P1, P2 => P2, Co => pout);

end SYN_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity PG_6 is

   port( G1, P1, G2, P2 : in std_logic;  gout, pout : out std_logic);

end PG_6;

architecture SYN_arch of PG_6 is

   component P_6
      port( p1, P2 : in std_logic;  Co : out std_logic);
   end component;
   
   component G_6
      port( G1, P, G2 : in std_logic;  Co : out std_logic);
   end component;

begin
   
   g_comp : G_6 port map( G1 => G1, P => P1, G2 => G2, Co => gout);
   p_comp : P_6 port map( p1 => P1, P2 => P2, Co => pout);

end SYN_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity PG_5 is

   port( G1, P1, G2, P2 : in std_logic;  gout, pout : out std_logic);

end PG_5;

architecture SYN_arch of PG_5 is

   component P_5
      port( p1, P2 : in std_logic;  Co : out std_logic);
   end component;
   
   component G_5
      port( G1, P, G2 : in std_logic;  Co : out std_logic);
   end component;

begin
   
   g_comp : G_5 port map( G1 => G1, P => P1, G2 => G2, Co => gout);
   p_comp : P_5 port map( p1 => P1, P2 => P2, Co => pout);

end SYN_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity PG_4 is

   port( G1, P1, G2, P2 : in std_logic;  gout, pout : out std_logic);

end PG_4;

architecture SYN_arch of PG_4 is

   component P_4
      port( p1, P2 : in std_logic;  Co : out std_logic);
   end component;
   
   component G_4
      port( G1, P, G2 : in std_logic;  Co : out std_logic);
   end component;

begin
   
   g_comp : G_4 port map( G1 => G1, P => P1, G2 => G2, Co => gout);
   p_comp : P_4 port map( p1 => P1, P2 => P2, Co => pout);

end SYN_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity PG_3 is

   port( G1, P1, G2, P2 : in std_logic;  gout, pout : out std_logic);

end PG_3;

architecture SYN_arch of PG_3 is

   component P_3
      port( p1, P2 : in std_logic;  Co : out std_logic);
   end component;
   
   component G_3
      port( G1, P, G2 : in std_logic;  Co : out std_logic);
   end component;

begin
   
   g_comp : G_3 port map( G1 => G1, P => P1, G2 => G2, Co => gout);
   p_comp : P_3 port map( p1 => P1, P2 => P2, Co => pout);

end SYN_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity PG_2 is

   port( G1, P1, G2, P2 : in std_logic;  gout, pout : out std_logic);

end PG_2;

architecture SYN_arch of PG_2 is

   component P_2
      port( p1, P2 : in std_logic;  Co : out std_logic);
   end component;
   
   component G_2
      port( G1, P, G2 : in std_logic;  Co : out std_logic);
   end component;

begin
   
   g_comp : G_2 port map( G1 => G1, P => P1, G2 => G2, Co => gout);
   p_comp : P_2 port map( p1 => P1, P2 => P2, Co => pout);

end SYN_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity PG_1 is

   port( G1, P1, G2, P2 : in std_logic;  gout, pout : out std_logic);

end PG_1;

architecture SYN_arch of PG_1 is

   component P_1
      port( p1, P2 : in std_logic;  Co : out std_logic);
   end component;
   
   component G_1
      port( G1, P, G2 : in std_logic;  Co : out std_logic);
   end component;

begin
   
   g_comp : G_1 port map( G1 => G1, P => P1, G2 => G2, Co => gout);
   p_comp : P_1 port map( p1 => P1, P2 => P2, Co => pout);

end SYN_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity G_52 is

   port( G1, P, G2 : in std_logic;  Co : out std_logic);

end G_52;

architecture SYN_behave of G_52 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => Co);
   U2 : AOI21_X1 port map( B1 => P, B2 => G2, A => G1, ZN => n3);

end SYN_behave;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity G_51 is

   port( G1, P, G2 : in std_logic;  Co : out std_logic);

end G_51;

architecture SYN_behave of G_51 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => Co);
   U2 : AOI21_X1 port map( B1 => P, B2 => G2, A => G1, ZN => n3);

end SYN_behave;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity G_50 is

   port( G1, P, G2 : in std_logic;  Co : out std_logic);

end G_50;

architecture SYN_behave of G_50 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => Co);
   U2 : AOI21_X1 port map( B1 => P, B2 => G2, A => G1, ZN => n3);

end SYN_behave;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity G_49 is

   port( G1, P, G2 : in std_logic;  Co : out std_logic);

end G_49;

architecture SYN_behave of G_49 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => Co);
   U2 : AOI21_X1 port map( B1 => P, B2 => G2, A => G1, ZN => n3);

end SYN_behave;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity G_48 is

   port( G1, P, G2 : in std_logic;  Co : out std_logic);

end G_48;

architecture SYN_behave of G_48 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => Co);
   U2 : AOI21_X1 port map( B1 => P, B2 => G2, A => G1, ZN => n3);

end SYN_behave;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity G_47 is

   port( G1, P, G2 : in std_logic;  Co : out std_logic);

end G_47;

architecture SYN_behave of G_47 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => Co);
   U2 : AOI21_X1 port map( B1 => P, B2 => G2, A => G1, ZN => n3);

end SYN_behave;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity G_46 is

   port( G1, P, G2 : in std_logic;  Co : out std_logic);

end G_46;

architecture SYN_behave of G_46 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => Co);
   U2 : AOI21_X1 port map( B1 => P, B2 => G2, A => G1, ZN => n3);

end SYN_behave;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity G_45 is

   port( G1, P, G2 : in std_logic;  Co : out std_logic);

end G_45;

architecture SYN_behave of G_45 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => Co);
   U2 : AOI21_X1 port map( B1 => P, B2 => G2, A => G1, ZN => n3);

end SYN_behave;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity G_44 is

   port( G1, P, G2 : in std_logic;  Co : out std_logic);

end G_44;

architecture SYN_behave of G_44 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => Co);
   U2 : AOI21_X1 port map( B1 => P, B2 => G2, A => G1, ZN => n3);

end SYN_behave;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity G_43 is

   port( G1, P, G2 : in std_logic;  Co : out std_logic);

end G_43;

architecture SYN_behave of G_43 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => Co);
   U2 : AOI21_X1 port map( B1 => P, B2 => G2, A => G1, ZN => n3);

end SYN_behave;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity G_42 is

   port( G1, P, G2 : in std_logic;  Co : out std_logic);

end G_42;

architecture SYN_behave of G_42 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => Co);
   U2 : AOI21_X1 port map( B1 => P, B2 => G2, A => G1, ZN => n3);

end SYN_behave;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity G_41 is

   port( G1, P, G2 : in std_logic;  Co : out std_logic);

end G_41;

architecture SYN_behave of G_41 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => Co);
   U2 : AOI21_X1 port map( B1 => P, B2 => G2, A => G1, ZN => n3);

end SYN_behave;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity G_40 is

   port( G1, P, G2 : in std_logic;  Co : out std_logic);

end G_40;

architecture SYN_behave of G_40 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => Co);
   U2 : AOI21_X1 port map( B1 => P, B2 => G2, A => G1, ZN => n3);

end SYN_behave;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity G_39 is

   port( G1, P, G2 : in std_logic;  Co : out std_logic);

end G_39;

architecture SYN_behave of G_39 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => Co);
   U2 : AOI21_X1 port map( B1 => P, B2 => G2, A => G1, ZN => n3);

end SYN_behave;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity G_38 is

   port( G1, P, G2 : in std_logic;  Co : out std_logic);

end G_38;

architecture SYN_behave of G_38 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => Co);
   U2 : AOI21_X1 port map( B1 => P, B2 => G2, A => G1, ZN => n3);

end SYN_behave;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity G_37 is

   port( G1, P, G2 : in std_logic;  Co : out std_logic);

end G_37;

architecture SYN_behave of G_37 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => Co);
   U2 : AOI21_X1 port map( B1 => P, B2 => G2, A => G1, ZN => n3);

end SYN_behave;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity G_36 is

   port( G1, P, G2 : in std_logic;  Co : out std_logic);

end G_36;

architecture SYN_behave of G_36 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => Co);
   U2 : AOI21_X1 port map( B1 => P, B2 => G2, A => G1, ZN => n3);

end SYN_behave;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity G_35 is

   port( G1, P, G2 : in std_logic;  Co : out std_logic);

end G_35;

architecture SYN_behave of G_35 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => Co);
   U2 : AOI21_X1 port map( B1 => P, B2 => G2, A => G1, ZN => n3);

end SYN_behave;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity G_34 is

   port( G1, P, G2 : in std_logic;  Co : out std_logic);

end G_34;

architecture SYN_behave of G_34 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => Co);
   U2 : AOI21_X1 port map( B1 => P, B2 => G2, A => G1, ZN => n3);

end SYN_behave;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity G_33 is

   port( G1, P, G2 : in std_logic;  Co : out std_logic);

end G_33;

architecture SYN_behave of G_33 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => Co);
   U2 : AOI21_X1 port map( B1 => P, B2 => G2, A => G1, ZN => n3);

end SYN_behave;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity G_32 is

   port( G1, P, G2 : in std_logic;  Co : out std_logic);

end G_32;

architecture SYN_behave of G_32 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => Co);
   U2 : AOI21_X1 port map( B1 => P, B2 => G2, A => G1, ZN => n3);

end SYN_behave;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity G_31 is

   port( G1, P, G2 : in std_logic;  Co : out std_logic);

end G_31;

architecture SYN_behave of G_31 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => Co);
   U2 : AOI21_X1 port map( B1 => P, B2 => G2, A => G1, ZN => n3);

end SYN_behave;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity G_30 is

   port( G1, P, G2 : in std_logic;  Co : out std_logic);

end G_30;

architecture SYN_behave of G_30 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => Co);
   U2 : AOI21_X1 port map( B1 => P, B2 => G2, A => G1, ZN => n3);

end SYN_behave;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity G_29 is

   port( G1, P, G2 : in std_logic;  Co : out std_logic);

end G_29;

architecture SYN_behave of G_29 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => Co);
   U2 : AOI21_X1 port map( B1 => P, B2 => G2, A => G1, ZN => n3);

end SYN_behave;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity G_28 is

   port( G1, P, G2 : in std_logic;  Co : out std_logic);

end G_28;

architecture SYN_behave of G_28 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => Co);
   U2 : AOI21_X1 port map( B1 => P, B2 => G2, A => G1, ZN => n3);

end SYN_behave;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity G_27 is

   port( G1, P, G2 : in std_logic;  Co : out std_logic);

end G_27;

architecture SYN_behave of G_27 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => Co);
   U2 : AOI21_X1 port map( B1 => P, B2 => G2, A => G1, ZN => n3);

end SYN_behave;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity G_26 is

   port( G1, P, G2 : in std_logic;  Co : out std_logic);

end G_26;

architecture SYN_behave of G_26 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => Co);
   U2 : AOI21_X1 port map( B1 => P, B2 => G2, A => G1, ZN => n3);

end SYN_behave;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity G_25 is

   port( G1, P, G2 : in std_logic;  Co : out std_logic);

end G_25;

architecture SYN_behave of G_25 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => Co);
   U2 : AOI21_X1 port map( B1 => P, B2 => G2, A => G1, ZN => n3);

end SYN_behave;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity G_24 is

   port( G1, P, G2 : in std_logic;  Co : out std_logic);

end G_24;

architecture SYN_behave of G_24 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => Co);
   U2 : AOI21_X1 port map( B1 => P, B2 => G2, A => G1, ZN => n3);

end SYN_behave;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity G_23 is

   port( G1, P, G2 : in std_logic;  Co : out std_logic);

end G_23;

architecture SYN_behave of G_23 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => Co);
   U2 : AOI21_X1 port map( B1 => P, B2 => G2, A => G1, ZN => n3);

end SYN_behave;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity G_22 is

   port( G1, P, G2 : in std_logic;  Co : out std_logic);

end G_22;

architecture SYN_behave of G_22 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => Co);
   U2 : AOI21_X1 port map( B1 => P, B2 => G2, A => G1, ZN => n3);

end SYN_behave;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity G_21 is

   port( G1, P, G2 : in std_logic;  Co : out std_logic);

end G_21;

architecture SYN_behave of G_21 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => Co);
   U2 : AOI21_X1 port map( B1 => P, B2 => G2, A => G1, ZN => n3);

end SYN_behave;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity G_20 is

   port( G1, P, G2 : in std_logic;  Co : out std_logic);

end G_20;

architecture SYN_behave of G_20 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => Co);
   U2 : AOI21_X1 port map( B1 => P, B2 => G2, A => G1, ZN => n3);

end SYN_behave;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity G_19 is

   port( G1, P, G2 : in std_logic;  Co : out std_logic);

end G_19;

architecture SYN_behave of G_19 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => Co);
   U2 : AOI21_X1 port map( B1 => P, B2 => G2, A => G1, ZN => n3);

end SYN_behave;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity G_18 is

   port( G1, P, G2 : in std_logic;  Co : out std_logic);

end G_18;

architecture SYN_behave of G_18 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => Co);
   U2 : AOI21_X1 port map( B1 => P, B2 => G2, A => G1, ZN => n3);

end SYN_behave;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity G_17 is

   port( G1, P, G2 : in std_logic;  Co : out std_logic);

end G_17;

architecture SYN_behave of G_17 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => Co);
   U2 : AOI21_X1 port map( B1 => P, B2 => G2, A => G1, ZN => n3);

end SYN_behave;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity G_16 is

   port( G1, P, G2 : in std_logic;  Co : out std_logic);

end G_16;

architecture SYN_behave of G_16 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => Co);
   U2 : AOI21_X1 port map( B1 => P, B2 => G2, A => G1, ZN => n3);

end SYN_behave;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity G_15 is

   port( G1, P, G2 : in std_logic;  Co : out std_logic);

end G_15;

architecture SYN_behave of G_15 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => Co);
   U2 : AOI21_X1 port map( B1 => P, B2 => G2, A => G1, ZN => n3);

end SYN_behave;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity G_14 is

   port( G1, P, G2 : in std_logic;  Co : out std_logic);

end G_14;

architecture SYN_behave of G_14 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => Co);
   U2 : AOI21_X1 port map( B1 => P, B2 => G2, A => G1, ZN => n3);

end SYN_behave;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity G_13 is

   port( G1, P, G2 : in std_logic;  Co : out std_logic);

end G_13;

architecture SYN_behave of G_13 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => Co);
   U2 : AOI21_X1 port map( B1 => P, B2 => G2, A => G1, ZN => n3);

end SYN_behave;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity G_12 is

   port( G1, P, G2 : in std_logic;  Co : out std_logic);

end G_12;

architecture SYN_behave of G_12 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => Co);
   U2 : AOI21_X1 port map( B1 => P, B2 => G2, A => G1, ZN => n3);

end SYN_behave;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity G_11 is

   port( G1, P, G2 : in std_logic;  Co : out std_logic);

end G_11;

architecture SYN_behave of G_11 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => Co);
   U2 : AOI21_X1 port map( B1 => P, B2 => G2, A => G1, ZN => n3);

end SYN_behave;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity G_10 is

   port( G1, P, G2 : in std_logic;  Co : out std_logic);

end G_10;

architecture SYN_behave of G_10 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => Co);
   U2 : AOI21_X1 port map( B1 => P, B2 => G2, A => G1, ZN => n3);

end SYN_behave;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity G_9 is

   port( G1, P, G2 : in std_logic;  Co : out std_logic);

end G_9;

architecture SYN_behave of G_9 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => Co);
   U2 : AOI21_X1 port map( B1 => P, B2 => G2, A => G1, ZN => n3);

end SYN_behave;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity G_8 is

   port( G1, P, G2 : in std_logic;  Co : out std_logic);

end G_8;

architecture SYN_behave of G_8 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => Co);
   U2 : AOI21_X1 port map( B1 => P, B2 => G2, A => G1, ZN => n3);

end SYN_behave;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity G_7 is

   port( G1, P, G2 : in std_logic;  Co : out std_logic);

end G_7;

architecture SYN_behave of G_7 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => Co);
   U2 : AOI21_X1 port map( B1 => P, B2 => G2, A => G1, ZN => n3);

end SYN_behave;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity G_6 is

   port( G1, P, G2 : in std_logic;  Co : out std_logic);

end G_6;

architecture SYN_behave of G_6 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => Co);
   U2 : AOI21_X1 port map( B1 => P, B2 => G2, A => G1, ZN => n3);

end SYN_behave;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity G_5 is

   port( G1, P, G2 : in std_logic;  Co : out std_logic);

end G_5;

architecture SYN_behave of G_5 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => Co);
   U2 : AOI21_X1 port map( B1 => P, B2 => G2, A => G1, ZN => n3);

end SYN_behave;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity G_4 is

   port( G1, P, G2 : in std_logic;  Co : out std_logic);

end G_4;

architecture SYN_behave of G_4 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => Co);
   U2 : AOI21_X1 port map( B1 => P, B2 => G2, A => G1, ZN => n3);

end SYN_behave;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity G_3 is

   port( G1, P, G2 : in std_logic;  Co : out std_logic);

end G_3;

architecture SYN_behave of G_3 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => Co);
   U2 : AOI21_X1 port map( B1 => P, B2 => G2, A => G1, ZN => n3);

end SYN_behave;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity G_2 is

   port( G1, P, G2 : in std_logic;  Co : out std_logic);

end G_2;

architecture SYN_behave of G_2 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => Co);
   U2 : AOI21_X1 port map( B1 => P, B2 => G2, A => G1, ZN => n3);

end SYN_behave;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity G_1 is

   port( G1, P, G2 : in std_logic;  Co : out std_logic);

end G_1;

architecture SYN_behave of G_1 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => Co);
   U2 : AOI21_X1 port map( B1 => P, B2 => G2, A => G1, ZN => n3);

end SYN_behave;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_767 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_767;

architecture SYN_ARCH2 of ND2_767 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_766 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_766;

architecture SYN_ARCH2 of ND2_766 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_765 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_765;

architecture SYN_ARCH2 of ND2_765 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_764 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_764;

architecture SYN_ARCH2 of ND2_764 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_763 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_763;

architecture SYN_ARCH2 of ND2_763 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_762 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_762;

architecture SYN_ARCH2 of ND2_762 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_761 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_761;

architecture SYN_ARCH2 of ND2_761 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_760 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_760;

architecture SYN_ARCH2 of ND2_760 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_759 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_759;

architecture SYN_ARCH2 of ND2_759 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_758 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_758;

architecture SYN_ARCH2 of ND2_758 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_757 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_757;

architecture SYN_ARCH2 of ND2_757 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_756 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_756;

architecture SYN_ARCH2 of ND2_756 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_755 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_755;

architecture SYN_ARCH2 of ND2_755 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_754 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_754;

architecture SYN_ARCH2 of ND2_754 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_753 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_753;

architecture SYN_ARCH2 of ND2_753 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_752 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_752;

architecture SYN_ARCH2 of ND2_752 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_751 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_751;

architecture SYN_ARCH2 of ND2_751 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_750 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_750;

architecture SYN_ARCH2 of ND2_750 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_749 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_749;

architecture SYN_ARCH2 of ND2_749 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_748 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_748;

architecture SYN_ARCH2 of ND2_748 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_747 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_747;

architecture SYN_ARCH2 of ND2_747 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_746 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_746;

architecture SYN_ARCH2 of ND2_746 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_745 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_745;

architecture SYN_ARCH2 of ND2_745 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_744 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_744;

architecture SYN_ARCH2 of ND2_744 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_743 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_743;

architecture SYN_ARCH2 of ND2_743 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_742 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_742;

architecture SYN_ARCH2 of ND2_742 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_741 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_741;

architecture SYN_ARCH2 of ND2_741 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_740 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_740;

architecture SYN_ARCH2 of ND2_740 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_739 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_739;

architecture SYN_ARCH2 of ND2_739 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_738 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_738;

architecture SYN_ARCH2 of ND2_738 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_737 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_737;

architecture SYN_ARCH2 of ND2_737 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_736 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_736;

architecture SYN_ARCH2 of ND2_736 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_735 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_735;

architecture SYN_ARCH2 of ND2_735 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_734 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_734;

architecture SYN_ARCH2 of ND2_734 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_733 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_733;

architecture SYN_ARCH2 of ND2_733 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_732 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_732;

architecture SYN_ARCH2 of ND2_732 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_731 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_731;

architecture SYN_ARCH2 of ND2_731 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_730 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_730;

architecture SYN_ARCH2 of ND2_730 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_729 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_729;

architecture SYN_ARCH2 of ND2_729 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_728 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_728;

architecture SYN_ARCH2 of ND2_728 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_727 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_727;

architecture SYN_ARCH2 of ND2_727 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_726 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_726;

architecture SYN_ARCH2 of ND2_726 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_725 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_725;

architecture SYN_ARCH2 of ND2_725 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_724 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_724;

architecture SYN_ARCH2 of ND2_724 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_723 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_723;

architecture SYN_ARCH2 of ND2_723 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_722 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_722;

architecture SYN_ARCH2 of ND2_722 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_721 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_721;

architecture SYN_ARCH2 of ND2_721 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_720 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_720;

architecture SYN_ARCH2 of ND2_720 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_719 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_719;

architecture SYN_ARCH2 of ND2_719 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_718 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_718;

architecture SYN_ARCH2 of ND2_718 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_717 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_717;

architecture SYN_ARCH2 of ND2_717 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_716 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_716;

architecture SYN_ARCH2 of ND2_716 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_715 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_715;

architecture SYN_ARCH2 of ND2_715 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_714 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_714;

architecture SYN_ARCH2 of ND2_714 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_713 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_713;

architecture SYN_ARCH2 of ND2_713 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_712 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_712;

architecture SYN_ARCH2 of ND2_712 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_711 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_711;

architecture SYN_ARCH2 of ND2_711 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_710 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_710;

architecture SYN_ARCH2 of ND2_710 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_709 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_709;

architecture SYN_ARCH2 of ND2_709 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_708 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_708;

architecture SYN_ARCH2 of ND2_708 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_707 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_707;

architecture SYN_ARCH2 of ND2_707 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_706 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_706;

architecture SYN_ARCH2 of ND2_706 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_705 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_705;

architecture SYN_ARCH2 of ND2_705 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_704 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_704;

architecture SYN_ARCH2 of ND2_704 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_703 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_703;

architecture SYN_ARCH2 of ND2_703 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_702 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_702;

architecture SYN_ARCH2 of ND2_702 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_701 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_701;

architecture SYN_ARCH2 of ND2_701 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_700 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_700;

architecture SYN_ARCH2 of ND2_700 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_699 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_699;

architecture SYN_ARCH2 of ND2_699 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_698 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_698;

architecture SYN_ARCH2 of ND2_698 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_697 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_697;

architecture SYN_ARCH2 of ND2_697 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_696 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_696;

architecture SYN_ARCH2 of ND2_696 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_695 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_695;

architecture SYN_ARCH2 of ND2_695 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_694 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_694;

architecture SYN_ARCH2 of ND2_694 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_693 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_693;

architecture SYN_ARCH2 of ND2_693 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_692 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_692;

architecture SYN_ARCH2 of ND2_692 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_691 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_691;

architecture SYN_ARCH2 of ND2_691 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_690 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_690;

architecture SYN_ARCH2 of ND2_690 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_689 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_689;

architecture SYN_ARCH2 of ND2_689 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_688 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_688;

architecture SYN_ARCH2 of ND2_688 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_687 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_687;

architecture SYN_ARCH2 of ND2_687 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_686 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_686;

architecture SYN_ARCH2 of ND2_686 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_685 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_685;

architecture SYN_ARCH2 of ND2_685 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_684 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_684;

architecture SYN_ARCH2 of ND2_684 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_683 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_683;

architecture SYN_ARCH2 of ND2_683 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_682 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_682;

architecture SYN_ARCH2 of ND2_682 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_681 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_681;

architecture SYN_ARCH2 of ND2_681 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_680 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_680;

architecture SYN_ARCH2 of ND2_680 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_679 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_679;

architecture SYN_ARCH2 of ND2_679 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_678 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_678;

architecture SYN_ARCH2 of ND2_678 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_677 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_677;

architecture SYN_ARCH2 of ND2_677 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_676 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_676;

architecture SYN_ARCH2 of ND2_676 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_675 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_675;

architecture SYN_ARCH2 of ND2_675 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_674 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_674;

architecture SYN_ARCH2 of ND2_674 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_673 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_673;

architecture SYN_ARCH2 of ND2_673 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_672 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_672;

architecture SYN_ARCH2 of ND2_672 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_671 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_671;

architecture SYN_ARCH2 of ND2_671 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_670 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_670;

architecture SYN_ARCH2 of ND2_670 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_669 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_669;

architecture SYN_ARCH2 of ND2_669 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_668 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_668;

architecture SYN_ARCH2 of ND2_668 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_667 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_667;

architecture SYN_ARCH2 of ND2_667 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_666 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_666;

architecture SYN_ARCH2 of ND2_666 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_665 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_665;

architecture SYN_ARCH2 of ND2_665 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_664 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_664;

architecture SYN_ARCH2 of ND2_664 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_663 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_663;

architecture SYN_ARCH2 of ND2_663 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_662 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_662;

architecture SYN_ARCH2 of ND2_662 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_661 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_661;

architecture SYN_ARCH2 of ND2_661 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_660 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_660;

architecture SYN_ARCH2 of ND2_660 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_659 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_659;

architecture SYN_ARCH2 of ND2_659 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_658 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_658;

architecture SYN_ARCH2 of ND2_658 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_657 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_657;

architecture SYN_ARCH2 of ND2_657 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_656 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_656;

architecture SYN_ARCH2 of ND2_656 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_655 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_655;

architecture SYN_ARCH2 of ND2_655 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_654 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_654;

architecture SYN_ARCH2 of ND2_654 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_653 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_653;

architecture SYN_ARCH2 of ND2_653 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_652 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_652;

architecture SYN_ARCH2 of ND2_652 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_651 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_651;

architecture SYN_ARCH2 of ND2_651 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_650 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_650;

architecture SYN_ARCH2 of ND2_650 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_649 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_649;

architecture SYN_ARCH2 of ND2_649 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_648 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_648;

architecture SYN_ARCH2 of ND2_648 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_647 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_647;

architecture SYN_ARCH2 of ND2_647 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_646 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_646;

architecture SYN_ARCH2 of ND2_646 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_645 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_645;

architecture SYN_ARCH2 of ND2_645 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_644 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_644;

architecture SYN_ARCH2 of ND2_644 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_643 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_643;

architecture SYN_ARCH2 of ND2_643 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_642 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_642;

architecture SYN_ARCH2 of ND2_642 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_641 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_641;

architecture SYN_ARCH2 of ND2_641 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_640 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_640;

architecture SYN_ARCH2 of ND2_640 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_639 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_639;

architecture SYN_ARCH2 of ND2_639 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_638 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_638;

architecture SYN_ARCH2 of ND2_638 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_637 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_637;

architecture SYN_ARCH2 of ND2_637 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_636 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_636;

architecture SYN_ARCH2 of ND2_636 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_635 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_635;

architecture SYN_ARCH2 of ND2_635 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_634 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_634;

architecture SYN_ARCH2 of ND2_634 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_633 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_633;

architecture SYN_ARCH2 of ND2_633 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_632 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_632;

architecture SYN_ARCH2 of ND2_632 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_631 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_631;

architecture SYN_ARCH2 of ND2_631 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_630 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_630;

architecture SYN_ARCH2 of ND2_630 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_629 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_629;

architecture SYN_ARCH2 of ND2_629 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_628 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_628;

architecture SYN_ARCH2 of ND2_628 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_627 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_627;

architecture SYN_ARCH2 of ND2_627 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_626 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_626;

architecture SYN_ARCH2 of ND2_626 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_625 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_625;

architecture SYN_ARCH2 of ND2_625 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_624 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_624;

architecture SYN_ARCH2 of ND2_624 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_623 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_623;

architecture SYN_ARCH2 of ND2_623 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_622 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_622;

architecture SYN_ARCH2 of ND2_622 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_621 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_621;

architecture SYN_ARCH2 of ND2_621 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_620 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_620;

architecture SYN_ARCH2 of ND2_620 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_619 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_619;

architecture SYN_ARCH2 of ND2_619 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_618 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_618;

architecture SYN_ARCH2 of ND2_618 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_617 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_617;

architecture SYN_ARCH2 of ND2_617 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_616 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_616;

architecture SYN_ARCH2 of ND2_616 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_615 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_615;

architecture SYN_ARCH2 of ND2_615 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_614 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_614;

architecture SYN_ARCH2 of ND2_614 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_613 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_613;

architecture SYN_ARCH2 of ND2_613 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_612 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_612;

architecture SYN_ARCH2 of ND2_612 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_611 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_611;

architecture SYN_ARCH2 of ND2_611 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_610 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_610;

architecture SYN_ARCH2 of ND2_610 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_609 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_609;

architecture SYN_ARCH2 of ND2_609 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_608 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_608;

architecture SYN_ARCH2 of ND2_608 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_607 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_607;

architecture SYN_ARCH2 of ND2_607 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_606 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_606;

architecture SYN_ARCH2 of ND2_606 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_605 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_605;

architecture SYN_ARCH2 of ND2_605 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_604 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_604;

architecture SYN_ARCH2 of ND2_604 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_603 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_603;

architecture SYN_ARCH2 of ND2_603 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_602 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_602;

architecture SYN_ARCH2 of ND2_602 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_601 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_601;

architecture SYN_ARCH2 of ND2_601 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_600 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_600;

architecture SYN_ARCH2 of ND2_600 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_599 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_599;

architecture SYN_ARCH2 of ND2_599 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_598 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_598;

architecture SYN_ARCH2 of ND2_598 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_597 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_597;

architecture SYN_ARCH2 of ND2_597 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_596 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_596;

architecture SYN_ARCH2 of ND2_596 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_595 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_595;

architecture SYN_ARCH2 of ND2_595 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_594 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_594;

architecture SYN_ARCH2 of ND2_594 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_593 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_593;

architecture SYN_ARCH2 of ND2_593 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_592 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_592;

architecture SYN_ARCH2 of ND2_592 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_591 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_591;

architecture SYN_ARCH2 of ND2_591 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_590 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_590;

architecture SYN_ARCH2 of ND2_590 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_589 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_589;

architecture SYN_ARCH2 of ND2_589 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_588 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_588;

architecture SYN_ARCH2 of ND2_588 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_587 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_587;

architecture SYN_ARCH2 of ND2_587 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_586 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_586;

architecture SYN_ARCH2 of ND2_586 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_585 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_585;

architecture SYN_ARCH2 of ND2_585 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_584 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_584;

architecture SYN_ARCH2 of ND2_584 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_583 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_583;

architecture SYN_ARCH2 of ND2_583 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_582 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_582;

architecture SYN_ARCH2 of ND2_582 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_581 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_581;

architecture SYN_ARCH2 of ND2_581 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_580 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_580;

architecture SYN_ARCH2 of ND2_580 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_579 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_579;

architecture SYN_ARCH2 of ND2_579 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_578 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_578;

architecture SYN_ARCH2 of ND2_578 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_577 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_577;

architecture SYN_ARCH2 of ND2_577 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_576 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_576;

architecture SYN_ARCH2 of ND2_576 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_575 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_575;

architecture SYN_ARCH2 of ND2_575 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_574 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_574;

architecture SYN_ARCH2 of ND2_574 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_573 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_573;

architecture SYN_ARCH2 of ND2_573 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_572 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_572;

architecture SYN_ARCH2 of ND2_572 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_571 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_571;

architecture SYN_ARCH2 of ND2_571 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_570 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_570;

architecture SYN_ARCH2 of ND2_570 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_569 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_569;

architecture SYN_ARCH2 of ND2_569 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_568 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_568;

architecture SYN_ARCH2 of ND2_568 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_567 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_567;

architecture SYN_ARCH2 of ND2_567 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_566 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_566;

architecture SYN_ARCH2 of ND2_566 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_565 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_565;

architecture SYN_ARCH2 of ND2_565 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_564 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_564;

architecture SYN_ARCH2 of ND2_564 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_563 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_563;

architecture SYN_ARCH2 of ND2_563 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_562 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_562;

architecture SYN_ARCH2 of ND2_562 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_561 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_561;

architecture SYN_ARCH2 of ND2_561 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_560 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_560;

architecture SYN_ARCH2 of ND2_560 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_559 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_559;

architecture SYN_ARCH2 of ND2_559 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_558 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_558;

architecture SYN_ARCH2 of ND2_558 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_557 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_557;

architecture SYN_ARCH2 of ND2_557 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_556 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_556;

architecture SYN_ARCH2 of ND2_556 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_555 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_555;

architecture SYN_ARCH2 of ND2_555 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_554 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_554;

architecture SYN_ARCH2 of ND2_554 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_553 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_553;

architecture SYN_ARCH2 of ND2_553 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_552 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_552;

architecture SYN_ARCH2 of ND2_552 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_551 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_551;

architecture SYN_ARCH2 of ND2_551 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_550 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_550;

architecture SYN_ARCH2 of ND2_550 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_549 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_549;

architecture SYN_ARCH2 of ND2_549 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_548 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_548;

architecture SYN_ARCH2 of ND2_548 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_547 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_547;

architecture SYN_ARCH2 of ND2_547 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_546 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_546;

architecture SYN_ARCH2 of ND2_546 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_545 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_545;

architecture SYN_ARCH2 of ND2_545 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_544 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_544;

architecture SYN_ARCH2 of ND2_544 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_543 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_543;

architecture SYN_ARCH2 of ND2_543 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_542 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_542;

architecture SYN_ARCH2 of ND2_542 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_541 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_541;

architecture SYN_ARCH2 of ND2_541 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_540 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_540;

architecture SYN_ARCH2 of ND2_540 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_539 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_539;

architecture SYN_ARCH2 of ND2_539 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_538 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_538;

architecture SYN_ARCH2 of ND2_538 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_537 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_537;

architecture SYN_ARCH2 of ND2_537 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_536 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_536;

architecture SYN_ARCH2 of ND2_536 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_535 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_535;

architecture SYN_ARCH2 of ND2_535 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_534 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_534;

architecture SYN_ARCH2 of ND2_534 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_533 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_533;

architecture SYN_ARCH2 of ND2_533 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_532 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_532;

architecture SYN_ARCH2 of ND2_532 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_531 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_531;

architecture SYN_ARCH2 of ND2_531 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_530 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_530;

architecture SYN_ARCH2 of ND2_530 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_529 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_529;

architecture SYN_ARCH2 of ND2_529 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_528 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_528;

architecture SYN_ARCH2 of ND2_528 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_527 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_527;

architecture SYN_ARCH2 of ND2_527 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_526 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_526;

architecture SYN_ARCH2 of ND2_526 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_525 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_525;

architecture SYN_ARCH2 of ND2_525 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_524 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_524;

architecture SYN_ARCH2 of ND2_524 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_523 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_523;

architecture SYN_ARCH2 of ND2_523 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_522 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_522;

architecture SYN_ARCH2 of ND2_522 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_521 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_521;

architecture SYN_ARCH2 of ND2_521 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_520 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_520;

architecture SYN_ARCH2 of ND2_520 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_519 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_519;

architecture SYN_ARCH2 of ND2_519 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_518 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_518;

architecture SYN_ARCH2 of ND2_518 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_517 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_517;

architecture SYN_ARCH2 of ND2_517 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_516 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_516;

architecture SYN_ARCH2 of ND2_516 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_515 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_515;

architecture SYN_ARCH2 of ND2_515 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_514 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_514;

architecture SYN_ARCH2 of ND2_514 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_513 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_513;

architecture SYN_ARCH2 of ND2_513 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_512 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_512;

architecture SYN_ARCH2 of ND2_512 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_511 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_511;

architecture SYN_ARCH2 of ND2_511 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_510 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_510;

architecture SYN_ARCH2 of ND2_510 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_509 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_509;

architecture SYN_ARCH2 of ND2_509 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_508 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_508;

architecture SYN_ARCH2 of ND2_508 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_507 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_507;

architecture SYN_ARCH2 of ND2_507 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_506 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_506;

architecture SYN_ARCH2 of ND2_506 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_505 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_505;

architecture SYN_ARCH2 of ND2_505 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_504 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_504;

architecture SYN_ARCH2 of ND2_504 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_503 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_503;

architecture SYN_ARCH2 of ND2_503 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_502 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_502;

architecture SYN_ARCH2 of ND2_502 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_501 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_501;

architecture SYN_ARCH2 of ND2_501 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_500 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_500;

architecture SYN_ARCH2 of ND2_500 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_499 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_499;

architecture SYN_ARCH2 of ND2_499 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_498 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_498;

architecture SYN_ARCH2 of ND2_498 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_497 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_497;

architecture SYN_ARCH2 of ND2_497 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_496 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_496;

architecture SYN_ARCH2 of ND2_496 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_495 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_495;

architecture SYN_ARCH2 of ND2_495 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_494 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_494;

architecture SYN_ARCH2 of ND2_494 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_493 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_493;

architecture SYN_ARCH2 of ND2_493 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_492 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_492;

architecture SYN_ARCH2 of ND2_492 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_491 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_491;

architecture SYN_ARCH2 of ND2_491 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_490 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_490;

architecture SYN_ARCH2 of ND2_490 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_489 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_489;

architecture SYN_ARCH2 of ND2_489 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_488 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_488;

architecture SYN_ARCH2 of ND2_488 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_487 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_487;

architecture SYN_ARCH2 of ND2_487 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_486 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_486;

architecture SYN_ARCH2 of ND2_486 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_485 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_485;

architecture SYN_ARCH2 of ND2_485 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_484 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_484;

architecture SYN_ARCH2 of ND2_484 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_483 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_483;

architecture SYN_ARCH2 of ND2_483 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_482 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_482;

architecture SYN_ARCH2 of ND2_482 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_481 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_481;

architecture SYN_ARCH2 of ND2_481 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_480 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_480;

architecture SYN_ARCH2 of ND2_480 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_479 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_479;

architecture SYN_ARCH2 of ND2_479 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_478 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_478;

architecture SYN_ARCH2 of ND2_478 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_477 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_477;

architecture SYN_ARCH2 of ND2_477 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_476 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_476;

architecture SYN_ARCH2 of ND2_476 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_475 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_475;

architecture SYN_ARCH2 of ND2_475 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_474 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_474;

architecture SYN_ARCH2 of ND2_474 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_473 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_473;

architecture SYN_ARCH2 of ND2_473 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_472 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_472;

architecture SYN_ARCH2 of ND2_472 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_471 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_471;

architecture SYN_ARCH2 of ND2_471 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_470 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_470;

architecture SYN_ARCH2 of ND2_470 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_469 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_469;

architecture SYN_ARCH2 of ND2_469 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_468 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_468;

architecture SYN_ARCH2 of ND2_468 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_467 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_467;

architecture SYN_ARCH2 of ND2_467 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_466 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_466;

architecture SYN_ARCH2 of ND2_466 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_465 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_465;

architecture SYN_ARCH2 of ND2_465 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_464 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_464;

architecture SYN_ARCH2 of ND2_464 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_463 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_463;

architecture SYN_ARCH2 of ND2_463 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_462 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_462;

architecture SYN_ARCH2 of ND2_462 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_461 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_461;

architecture SYN_ARCH2 of ND2_461 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_460 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_460;

architecture SYN_ARCH2 of ND2_460 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_459 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_459;

architecture SYN_ARCH2 of ND2_459 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_458 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_458;

architecture SYN_ARCH2 of ND2_458 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_457 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_457;

architecture SYN_ARCH2 of ND2_457 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_456 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_456;

architecture SYN_ARCH2 of ND2_456 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_455 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_455;

architecture SYN_ARCH2 of ND2_455 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_454 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_454;

architecture SYN_ARCH2 of ND2_454 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_453 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_453;

architecture SYN_ARCH2 of ND2_453 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_452 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_452;

architecture SYN_ARCH2 of ND2_452 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_451 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_451;

architecture SYN_ARCH2 of ND2_451 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_450 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_450;

architecture SYN_ARCH2 of ND2_450 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_449 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_449;

architecture SYN_ARCH2 of ND2_449 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_448 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_448;

architecture SYN_ARCH2 of ND2_448 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_447 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_447;

architecture SYN_ARCH2 of ND2_447 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_446 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_446;

architecture SYN_ARCH2 of ND2_446 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_445 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_445;

architecture SYN_ARCH2 of ND2_445 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_444 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_444;

architecture SYN_ARCH2 of ND2_444 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_443 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_443;

architecture SYN_ARCH2 of ND2_443 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_442 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_442;

architecture SYN_ARCH2 of ND2_442 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_441 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_441;

architecture SYN_ARCH2 of ND2_441 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_440 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_440;

architecture SYN_ARCH2 of ND2_440 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_439 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_439;

architecture SYN_ARCH2 of ND2_439 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_438 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_438;

architecture SYN_ARCH2 of ND2_438 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_437 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_437;

architecture SYN_ARCH2 of ND2_437 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_436 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_436;

architecture SYN_ARCH2 of ND2_436 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_435 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_435;

architecture SYN_ARCH2 of ND2_435 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_434 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_434;

architecture SYN_ARCH2 of ND2_434 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_433 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_433;

architecture SYN_ARCH2 of ND2_433 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_432 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_432;

architecture SYN_ARCH2 of ND2_432 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_431 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_431;

architecture SYN_ARCH2 of ND2_431 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_430 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_430;

architecture SYN_ARCH2 of ND2_430 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_429 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_429;

architecture SYN_ARCH2 of ND2_429 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_428 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_428;

architecture SYN_ARCH2 of ND2_428 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_427 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_427;

architecture SYN_ARCH2 of ND2_427 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_426 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_426;

architecture SYN_ARCH2 of ND2_426 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_425 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_425;

architecture SYN_ARCH2 of ND2_425 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_424 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_424;

architecture SYN_ARCH2 of ND2_424 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_423 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_423;

architecture SYN_ARCH2 of ND2_423 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_422 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_422;

architecture SYN_ARCH2 of ND2_422 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_421 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_421;

architecture SYN_ARCH2 of ND2_421 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_420 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_420;

architecture SYN_ARCH2 of ND2_420 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_419 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_419;

architecture SYN_ARCH2 of ND2_419 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_418 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_418;

architecture SYN_ARCH2 of ND2_418 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_417 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_417;

architecture SYN_ARCH2 of ND2_417 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_416 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_416;

architecture SYN_ARCH2 of ND2_416 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_415 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_415;

architecture SYN_ARCH2 of ND2_415 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_414 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_414;

architecture SYN_ARCH2 of ND2_414 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_413 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_413;

architecture SYN_ARCH2 of ND2_413 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_412 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_412;

architecture SYN_ARCH2 of ND2_412 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_411 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_411;

architecture SYN_ARCH2 of ND2_411 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_410 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_410;

architecture SYN_ARCH2 of ND2_410 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_409 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_409;

architecture SYN_ARCH2 of ND2_409 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_408 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_408;

architecture SYN_ARCH2 of ND2_408 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_407 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_407;

architecture SYN_ARCH2 of ND2_407 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_406 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_406;

architecture SYN_ARCH2 of ND2_406 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_405 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_405;

architecture SYN_ARCH2 of ND2_405 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_404 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_404;

architecture SYN_ARCH2 of ND2_404 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_403 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_403;

architecture SYN_ARCH2 of ND2_403 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_402 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_402;

architecture SYN_ARCH2 of ND2_402 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_401 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_401;

architecture SYN_ARCH2 of ND2_401 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_400 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_400;

architecture SYN_ARCH2 of ND2_400 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_399 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_399;

architecture SYN_ARCH2 of ND2_399 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_398 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_398;

architecture SYN_ARCH2 of ND2_398 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_397 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_397;

architecture SYN_ARCH2 of ND2_397 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_396 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_396;

architecture SYN_ARCH2 of ND2_396 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_395 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_395;

architecture SYN_ARCH2 of ND2_395 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_394 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_394;

architecture SYN_ARCH2 of ND2_394 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_393 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_393;

architecture SYN_ARCH2 of ND2_393 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_392 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_392;

architecture SYN_ARCH2 of ND2_392 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_391 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_391;

architecture SYN_ARCH2 of ND2_391 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_390 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_390;

architecture SYN_ARCH2 of ND2_390 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_389 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_389;

architecture SYN_ARCH2 of ND2_389 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_388 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_388;

architecture SYN_ARCH2 of ND2_388 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_387 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_387;

architecture SYN_ARCH2 of ND2_387 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_386 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_386;

architecture SYN_ARCH2 of ND2_386 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_385 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_385;

architecture SYN_ARCH2 of ND2_385 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_384 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_384;

architecture SYN_ARCH2 of ND2_384 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_383 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_383;

architecture SYN_ARCH2 of ND2_383 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_382 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_382;

architecture SYN_ARCH2 of ND2_382 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_381 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_381;

architecture SYN_ARCH2 of ND2_381 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_380 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_380;

architecture SYN_ARCH2 of ND2_380 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_379 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_379;

architecture SYN_ARCH2 of ND2_379 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_378 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_378;

architecture SYN_ARCH2 of ND2_378 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_377 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_377;

architecture SYN_ARCH2 of ND2_377 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_376 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_376;

architecture SYN_ARCH2 of ND2_376 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_375 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_375;

architecture SYN_ARCH2 of ND2_375 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_374 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_374;

architecture SYN_ARCH2 of ND2_374 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_373 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_373;

architecture SYN_ARCH2 of ND2_373 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_372 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_372;

architecture SYN_ARCH2 of ND2_372 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_371 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_371;

architecture SYN_ARCH2 of ND2_371 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_370 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_370;

architecture SYN_ARCH2 of ND2_370 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_369 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_369;

architecture SYN_ARCH2 of ND2_369 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_368 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_368;

architecture SYN_ARCH2 of ND2_368 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_367 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_367;

architecture SYN_ARCH2 of ND2_367 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_366 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_366;

architecture SYN_ARCH2 of ND2_366 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_365 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_365;

architecture SYN_ARCH2 of ND2_365 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_364 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_364;

architecture SYN_ARCH2 of ND2_364 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_363 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_363;

architecture SYN_ARCH2 of ND2_363 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_362 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_362;

architecture SYN_ARCH2 of ND2_362 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_361 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_361;

architecture SYN_ARCH2 of ND2_361 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_360 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_360;

architecture SYN_ARCH2 of ND2_360 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_359 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_359;

architecture SYN_ARCH2 of ND2_359 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_358 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_358;

architecture SYN_ARCH2 of ND2_358 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_357 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_357;

architecture SYN_ARCH2 of ND2_357 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_356 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_356;

architecture SYN_ARCH2 of ND2_356 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_355 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_355;

architecture SYN_ARCH2 of ND2_355 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_354 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_354;

architecture SYN_ARCH2 of ND2_354 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_353 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_353;

architecture SYN_ARCH2 of ND2_353 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_352 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_352;

architecture SYN_ARCH2 of ND2_352 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_351 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_351;

architecture SYN_ARCH2 of ND2_351 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_350 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_350;

architecture SYN_ARCH2 of ND2_350 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_349 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_349;

architecture SYN_ARCH2 of ND2_349 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_348 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_348;

architecture SYN_ARCH2 of ND2_348 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_347 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_347;

architecture SYN_ARCH2 of ND2_347 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_346 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_346;

architecture SYN_ARCH2 of ND2_346 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_345 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_345;

architecture SYN_ARCH2 of ND2_345 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_344 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_344;

architecture SYN_ARCH2 of ND2_344 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_343 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_343;

architecture SYN_ARCH2 of ND2_343 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_342 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_342;

architecture SYN_ARCH2 of ND2_342 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_341 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_341;

architecture SYN_ARCH2 of ND2_341 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_340 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_340;

architecture SYN_ARCH2 of ND2_340 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_339 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_339;

architecture SYN_ARCH2 of ND2_339 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_338 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_338;

architecture SYN_ARCH2 of ND2_338 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_337 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_337;

architecture SYN_ARCH2 of ND2_337 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_336 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_336;

architecture SYN_ARCH2 of ND2_336 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_335 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_335;

architecture SYN_ARCH2 of ND2_335 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_334 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_334;

architecture SYN_ARCH2 of ND2_334 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_333 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_333;

architecture SYN_ARCH2 of ND2_333 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_332 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_332;

architecture SYN_ARCH2 of ND2_332 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_331 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_331;

architecture SYN_ARCH2 of ND2_331 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_330 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_330;

architecture SYN_ARCH2 of ND2_330 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_329 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_329;

architecture SYN_ARCH2 of ND2_329 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_328 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_328;

architecture SYN_ARCH2 of ND2_328 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_327 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_327;

architecture SYN_ARCH2 of ND2_327 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_326 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_326;

architecture SYN_ARCH2 of ND2_326 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_325 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_325;

architecture SYN_ARCH2 of ND2_325 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_324 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_324;

architecture SYN_ARCH2 of ND2_324 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_323 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_323;

architecture SYN_ARCH2 of ND2_323 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_322 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_322;

architecture SYN_ARCH2 of ND2_322 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_321 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_321;

architecture SYN_ARCH2 of ND2_321 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_320 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_320;

architecture SYN_ARCH2 of ND2_320 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_319 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_319;

architecture SYN_ARCH2 of ND2_319 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_318 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_318;

architecture SYN_ARCH2 of ND2_318 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_317 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_317;

architecture SYN_ARCH2 of ND2_317 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_316 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_316;

architecture SYN_ARCH2 of ND2_316 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_315 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_315;

architecture SYN_ARCH2 of ND2_315 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_314 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_314;

architecture SYN_ARCH2 of ND2_314 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_313 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_313;

architecture SYN_ARCH2 of ND2_313 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_312 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_312;

architecture SYN_ARCH2 of ND2_312 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_311 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_311;

architecture SYN_ARCH2 of ND2_311 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_310 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_310;

architecture SYN_ARCH2 of ND2_310 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_309 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_309;

architecture SYN_ARCH2 of ND2_309 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_308 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_308;

architecture SYN_ARCH2 of ND2_308 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_307 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_307;

architecture SYN_ARCH2 of ND2_307 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_306 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_306;

architecture SYN_ARCH2 of ND2_306 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_305 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_305;

architecture SYN_ARCH2 of ND2_305 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_304 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_304;

architecture SYN_ARCH2 of ND2_304 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_303 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_303;

architecture SYN_ARCH2 of ND2_303 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_302 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_302;

architecture SYN_ARCH2 of ND2_302 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_301 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_301;

architecture SYN_ARCH2 of ND2_301 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_300 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_300;

architecture SYN_ARCH2 of ND2_300 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_299 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_299;

architecture SYN_ARCH2 of ND2_299 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_298 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_298;

architecture SYN_ARCH2 of ND2_298 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_297 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_297;

architecture SYN_ARCH2 of ND2_297 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_296 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_296;

architecture SYN_ARCH2 of ND2_296 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_295 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_295;

architecture SYN_ARCH2 of ND2_295 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_294 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_294;

architecture SYN_ARCH2 of ND2_294 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_293 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_293;

architecture SYN_ARCH2 of ND2_293 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_292 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_292;

architecture SYN_ARCH2 of ND2_292 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_291 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_291;

architecture SYN_ARCH2 of ND2_291 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_290 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_290;

architecture SYN_ARCH2 of ND2_290 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_289 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_289;

architecture SYN_ARCH2 of ND2_289 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_288 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_288;

architecture SYN_ARCH2 of ND2_288 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_287 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_287;

architecture SYN_ARCH2 of ND2_287 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_286 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_286;

architecture SYN_ARCH2 of ND2_286 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_285 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_285;

architecture SYN_ARCH2 of ND2_285 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_284 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_284;

architecture SYN_ARCH2 of ND2_284 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_283 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_283;

architecture SYN_ARCH2 of ND2_283 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_282 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_282;

architecture SYN_ARCH2 of ND2_282 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_281 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_281;

architecture SYN_ARCH2 of ND2_281 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_280 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_280;

architecture SYN_ARCH2 of ND2_280 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_279 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_279;

architecture SYN_ARCH2 of ND2_279 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_278 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_278;

architecture SYN_ARCH2 of ND2_278 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_277 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_277;

architecture SYN_ARCH2 of ND2_277 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_276 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_276;

architecture SYN_ARCH2 of ND2_276 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_275 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_275;

architecture SYN_ARCH2 of ND2_275 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_274 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_274;

architecture SYN_ARCH2 of ND2_274 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_273 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_273;

architecture SYN_ARCH2 of ND2_273 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_272 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_272;

architecture SYN_ARCH2 of ND2_272 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_271 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_271;

architecture SYN_ARCH2 of ND2_271 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_270 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_270;

architecture SYN_ARCH2 of ND2_270 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_269 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_269;

architecture SYN_ARCH2 of ND2_269 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_268 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_268;

architecture SYN_ARCH2 of ND2_268 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_267 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_267;

architecture SYN_ARCH2 of ND2_267 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_266 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_266;

architecture SYN_ARCH2 of ND2_266 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_265 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_265;

architecture SYN_ARCH2 of ND2_265 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_264 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_264;

architecture SYN_ARCH2 of ND2_264 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_263 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_263;

architecture SYN_ARCH2 of ND2_263 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_262 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_262;

architecture SYN_ARCH2 of ND2_262 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_261 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_261;

architecture SYN_ARCH2 of ND2_261 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_260 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_260;

architecture SYN_ARCH2 of ND2_260 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_259 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_259;

architecture SYN_ARCH2 of ND2_259 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_258 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_258;

architecture SYN_ARCH2 of ND2_258 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_257 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_257;

architecture SYN_ARCH2 of ND2_257 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_256 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_256;

architecture SYN_ARCH2 of ND2_256 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_255 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_255;

architecture SYN_ARCH2 of ND2_255 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_254 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_254;

architecture SYN_ARCH2 of ND2_254 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_253 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_253;

architecture SYN_ARCH2 of ND2_253 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_252 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_252;

architecture SYN_ARCH2 of ND2_252 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_251 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_251;

architecture SYN_ARCH2 of ND2_251 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_250 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_250;

architecture SYN_ARCH2 of ND2_250 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_249 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_249;

architecture SYN_ARCH2 of ND2_249 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_248 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_248;

architecture SYN_ARCH2 of ND2_248 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_247 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_247;

architecture SYN_ARCH2 of ND2_247 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_246 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_246;

architecture SYN_ARCH2 of ND2_246 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_245 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_245;

architecture SYN_ARCH2 of ND2_245 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_244 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_244;

architecture SYN_ARCH2 of ND2_244 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_243 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_243;

architecture SYN_ARCH2 of ND2_243 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_242 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_242;

architecture SYN_ARCH2 of ND2_242 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_241 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_241;

architecture SYN_ARCH2 of ND2_241 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_240 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_240;

architecture SYN_ARCH2 of ND2_240 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_239 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_239;

architecture SYN_ARCH2 of ND2_239 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_238 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_238;

architecture SYN_ARCH2 of ND2_238 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_237 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_237;

architecture SYN_ARCH2 of ND2_237 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_236 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_236;

architecture SYN_ARCH2 of ND2_236 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_235 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_235;

architecture SYN_ARCH2 of ND2_235 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_234 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_234;

architecture SYN_ARCH2 of ND2_234 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_233 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_233;

architecture SYN_ARCH2 of ND2_233 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_232 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_232;

architecture SYN_ARCH2 of ND2_232 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_231 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_231;

architecture SYN_ARCH2 of ND2_231 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_230 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_230;

architecture SYN_ARCH2 of ND2_230 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_229 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_229;

architecture SYN_ARCH2 of ND2_229 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_228 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_228;

architecture SYN_ARCH2 of ND2_228 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_227 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_227;

architecture SYN_ARCH2 of ND2_227 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_226 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_226;

architecture SYN_ARCH2 of ND2_226 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_225 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_225;

architecture SYN_ARCH2 of ND2_225 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_224 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_224;

architecture SYN_ARCH2 of ND2_224 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_223 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_223;

architecture SYN_ARCH2 of ND2_223 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_222 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_222;

architecture SYN_ARCH2 of ND2_222 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_221 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_221;

architecture SYN_ARCH2 of ND2_221 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_220 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_220;

architecture SYN_ARCH2 of ND2_220 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_219 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_219;

architecture SYN_ARCH2 of ND2_219 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_218 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_218;

architecture SYN_ARCH2 of ND2_218 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_217 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_217;

architecture SYN_ARCH2 of ND2_217 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_216 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_216;

architecture SYN_ARCH2 of ND2_216 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_215 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_215;

architecture SYN_ARCH2 of ND2_215 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_214 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_214;

architecture SYN_ARCH2 of ND2_214 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_213 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_213;

architecture SYN_ARCH2 of ND2_213 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_212 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_212;

architecture SYN_ARCH2 of ND2_212 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_211 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_211;

architecture SYN_ARCH2 of ND2_211 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_210 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_210;

architecture SYN_ARCH2 of ND2_210 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_209 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_209;

architecture SYN_ARCH2 of ND2_209 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_208 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_208;

architecture SYN_ARCH2 of ND2_208 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_207 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_207;

architecture SYN_ARCH2 of ND2_207 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_206 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_206;

architecture SYN_ARCH2 of ND2_206 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_205 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_205;

architecture SYN_ARCH2 of ND2_205 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_204 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_204;

architecture SYN_ARCH2 of ND2_204 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_203 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_203;

architecture SYN_ARCH2 of ND2_203 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_202 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_202;

architecture SYN_ARCH2 of ND2_202 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_201 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_201;

architecture SYN_ARCH2 of ND2_201 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_200 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_200;

architecture SYN_ARCH2 of ND2_200 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_199 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_199;

architecture SYN_ARCH2 of ND2_199 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_198 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_198;

architecture SYN_ARCH2 of ND2_198 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_197 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_197;

architecture SYN_ARCH2 of ND2_197 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_196 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_196;

architecture SYN_ARCH2 of ND2_196 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_195 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_195;

architecture SYN_ARCH2 of ND2_195 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_194 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_194;

architecture SYN_ARCH2 of ND2_194 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_193 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_193;

architecture SYN_ARCH2 of ND2_193 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_192 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_192;

architecture SYN_ARCH2 of ND2_192 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_191 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_191;

architecture SYN_ARCH2 of ND2_191 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_190 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_190;

architecture SYN_ARCH2 of ND2_190 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_189 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_189;

architecture SYN_ARCH2 of ND2_189 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_188 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_188;

architecture SYN_ARCH2 of ND2_188 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_187 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_187;

architecture SYN_ARCH2 of ND2_187 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_186 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_186;

architecture SYN_ARCH2 of ND2_186 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_185 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_185;

architecture SYN_ARCH2 of ND2_185 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_184 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_184;

architecture SYN_ARCH2 of ND2_184 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_183 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_183;

architecture SYN_ARCH2 of ND2_183 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_182 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_182;

architecture SYN_ARCH2 of ND2_182 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_181 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_181;

architecture SYN_ARCH2 of ND2_181 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_180 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_180;

architecture SYN_ARCH2 of ND2_180 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_179 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_179;

architecture SYN_ARCH2 of ND2_179 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_178 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_178;

architecture SYN_ARCH2 of ND2_178 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_177 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_177;

architecture SYN_ARCH2 of ND2_177 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_176 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_176;

architecture SYN_ARCH2 of ND2_176 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_175 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_175;

architecture SYN_ARCH2 of ND2_175 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_174 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_174;

architecture SYN_ARCH2 of ND2_174 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_173 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_173;

architecture SYN_ARCH2 of ND2_173 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_172 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_172;

architecture SYN_ARCH2 of ND2_172 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_171 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_171;

architecture SYN_ARCH2 of ND2_171 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_170 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_170;

architecture SYN_ARCH2 of ND2_170 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_169 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_169;

architecture SYN_ARCH2 of ND2_169 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_168 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_168;

architecture SYN_ARCH2 of ND2_168 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_167 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_167;

architecture SYN_ARCH2 of ND2_167 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_166 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_166;

architecture SYN_ARCH2 of ND2_166 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_165 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_165;

architecture SYN_ARCH2 of ND2_165 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_164 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_164;

architecture SYN_ARCH2 of ND2_164 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_163 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_163;

architecture SYN_ARCH2 of ND2_163 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_162 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_162;

architecture SYN_ARCH2 of ND2_162 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_161 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_161;

architecture SYN_ARCH2 of ND2_161 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_160 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_160;

architecture SYN_ARCH2 of ND2_160 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_159 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_159;

architecture SYN_ARCH2 of ND2_159 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_158 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_158;

architecture SYN_ARCH2 of ND2_158 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_157 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_157;

architecture SYN_ARCH2 of ND2_157 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_156 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_156;

architecture SYN_ARCH2 of ND2_156 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_155 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_155;

architecture SYN_ARCH2 of ND2_155 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_154 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_154;

architecture SYN_ARCH2 of ND2_154 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_153 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_153;

architecture SYN_ARCH2 of ND2_153 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_152 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_152;

architecture SYN_ARCH2 of ND2_152 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_151 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_151;

architecture SYN_ARCH2 of ND2_151 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_150 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_150;

architecture SYN_ARCH2 of ND2_150 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_149 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_149;

architecture SYN_ARCH2 of ND2_149 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_148 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_148;

architecture SYN_ARCH2 of ND2_148 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_147 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_147;

architecture SYN_ARCH2 of ND2_147 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_146 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_146;

architecture SYN_ARCH2 of ND2_146 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_145 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_145;

architecture SYN_ARCH2 of ND2_145 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_144 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_144;

architecture SYN_ARCH2 of ND2_144 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_143 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_143;

architecture SYN_ARCH2 of ND2_143 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_142 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_142;

architecture SYN_ARCH2 of ND2_142 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_141 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_141;

architecture SYN_ARCH2 of ND2_141 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_140 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_140;

architecture SYN_ARCH2 of ND2_140 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_139 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_139;

architecture SYN_ARCH2 of ND2_139 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_138 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_138;

architecture SYN_ARCH2 of ND2_138 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_137 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_137;

architecture SYN_ARCH2 of ND2_137 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_136 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_136;

architecture SYN_ARCH2 of ND2_136 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_135 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_135;

architecture SYN_ARCH2 of ND2_135 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_134 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_134;

architecture SYN_ARCH2 of ND2_134 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_133 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_133;

architecture SYN_ARCH2 of ND2_133 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_132 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_132;

architecture SYN_ARCH2 of ND2_132 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_131 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_131;

architecture SYN_ARCH2 of ND2_131 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_130 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_130;

architecture SYN_ARCH2 of ND2_130 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_129 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_129;

architecture SYN_ARCH2 of ND2_129 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_128 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_128;

architecture SYN_ARCH2 of ND2_128 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_127 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_127;

architecture SYN_ARCH2 of ND2_127 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_126 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_126;

architecture SYN_ARCH2 of ND2_126 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_125 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_125;

architecture SYN_ARCH2 of ND2_125 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_124 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_124;

architecture SYN_ARCH2 of ND2_124 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_123 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_123;

architecture SYN_ARCH2 of ND2_123 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_122 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_122;

architecture SYN_ARCH2 of ND2_122 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_121 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_121;

architecture SYN_ARCH2 of ND2_121 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_120 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_120;

architecture SYN_ARCH2 of ND2_120 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_119 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_119;

architecture SYN_ARCH2 of ND2_119 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_118 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_118;

architecture SYN_ARCH2 of ND2_118 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_117 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_117;

architecture SYN_ARCH2 of ND2_117 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_116 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_116;

architecture SYN_ARCH2 of ND2_116 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_115 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_115;

architecture SYN_ARCH2 of ND2_115 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_114 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_114;

architecture SYN_ARCH2 of ND2_114 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_113 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_113;

architecture SYN_ARCH2 of ND2_113 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_112 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_112;

architecture SYN_ARCH2 of ND2_112 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_111 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_111;

architecture SYN_ARCH2 of ND2_111 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_110 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_110;

architecture SYN_ARCH2 of ND2_110 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_109 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_109;

architecture SYN_ARCH2 of ND2_109 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_108 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_108;

architecture SYN_ARCH2 of ND2_108 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_107 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_107;

architecture SYN_ARCH2 of ND2_107 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_106 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_106;

architecture SYN_ARCH2 of ND2_106 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_105 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_105;

architecture SYN_ARCH2 of ND2_105 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_104 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_104;

architecture SYN_ARCH2 of ND2_104 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_103 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_103;

architecture SYN_ARCH2 of ND2_103 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_102 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_102;

architecture SYN_ARCH2 of ND2_102 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_101 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_101;

architecture SYN_ARCH2 of ND2_101 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_100 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_100;

architecture SYN_ARCH2 of ND2_100 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_99 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_99;

architecture SYN_ARCH2 of ND2_99 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_98 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_98;

architecture SYN_ARCH2 of ND2_98 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_97 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_97;

architecture SYN_ARCH2 of ND2_97 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_96 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_96;

architecture SYN_ARCH2 of ND2_96 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_95 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_95;

architecture SYN_ARCH2 of ND2_95 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_94 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_94;

architecture SYN_ARCH2 of ND2_94 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_93 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_93;

architecture SYN_ARCH2 of ND2_93 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_92 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_92;

architecture SYN_ARCH2 of ND2_92 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_91 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_91;

architecture SYN_ARCH2 of ND2_91 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_90 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_90;

architecture SYN_ARCH2 of ND2_90 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_89 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_89;

architecture SYN_ARCH2 of ND2_89 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_88 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_88;

architecture SYN_ARCH2 of ND2_88 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_87 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_87;

architecture SYN_ARCH2 of ND2_87 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_86 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_86;

architecture SYN_ARCH2 of ND2_86 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_85 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_85;

architecture SYN_ARCH2 of ND2_85 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_84 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_84;

architecture SYN_ARCH2 of ND2_84 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_83 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_83;

architecture SYN_ARCH2 of ND2_83 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_82 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_82;

architecture SYN_ARCH2 of ND2_82 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_81 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_81;

architecture SYN_ARCH2 of ND2_81 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_80 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_80;

architecture SYN_ARCH2 of ND2_80 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_79 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_79;

architecture SYN_ARCH2 of ND2_79 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_78 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_78;

architecture SYN_ARCH2 of ND2_78 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_77 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_77;

architecture SYN_ARCH2 of ND2_77 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_76 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_76;

architecture SYN_ARCH2 of ND2_76 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_75 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_75;

architecture SYN_ARCH2 of ND2_75 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_74 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_74;

architecture SYN_ARCH2 of ND2_74 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_73 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_73;

architecture SYN_ARCH2 of ND2_73 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_72 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_72;

architecture SYN_ARCH2 of ND2_72 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_71 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_71;

architecture SYN_ARCH2 of ND2_71 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_70 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_70;

architecture SYN_ARCH2 of ND2_70 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_69 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_69;

architecture SYN_ARCH2 of ND2_69 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_68 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_68;

architecture SYN_ARCH2 of ND2_68 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_67 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_67;

architecture SYN_ARCH2 of ND2_67 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_66 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_66;

architecture SYN_ARCH2 of ND2_66 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_65 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_65;

architecture SYN_ARCH2 of ND2_65 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_64 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_64;

architecture SYN_ARCH2 of ND2_64 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_63 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_63;

architecture SYN_ARCH2 of ND2_63 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_62 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_62;

architecture SYN_ARCH2 of ND2_62 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_61 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_61;

architecture SYN_ARCH2 of ND2_61 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_60 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_60;

architecture SYN_ARCH2 of ND2_60 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_59 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_59;

architecture SYN_ARCH2 of ND2_59 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_58 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_58;

architecture SYN_ARCH2 of ND2_58 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_57 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_57;

architecture SYN_ARCH2 of ND2_57 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_56 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_56;

architecture SYN_ARCH2 of ND2_56 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_55 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_55;

architecture SYN_ARCH2 of ND2_55 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_54 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_54;

architecture SYN_ARCH2 of ND2_54 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_53 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_53;

architecture SYN_ARCH2 of ND2_53 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_52 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_52;

architecture SYN_ARCH2 of ND2_52 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_51 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_51;

architecture SYN_ARCH2 of ND2_51 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_50 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_50;

architecture SYN_ARCH2 of ND2_50 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_49 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_49;

architecture SYN_ARCH2 of ND2_49 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_48 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_48;

architecture SYN_ARCH2 of ND2_48 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_47 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_47;

architecture SYN_ARCH2 of ND2_47 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_46 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_46;

architecture SYN_ARCH2 of ND2_46 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_45 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_45;

architecture SYN_ARCH2 of ND2_45 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_44 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_44;

architecture SYN_ARCH2 of ND2_44 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_43 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_43;

architecture SYN_ARCH2 of ND2_43 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_42 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_42;

architecture SYN_ARCH2 of ND2_42 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_41 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_41;

architecture SYN_ARCH2 of ND2_41 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_40 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_40;

architecture SYN_ARCH2 of ND2_40 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_39 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_39;

architecture SYN_ARCH2 of ND2_39 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_38 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_38;

architecture SYN_ARCH2 of ND2_38 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_37 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_37;

architecture SYN_ARCH2 of ND2_37 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_36 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_36;

architecture SYN_ARCH2 of ND2_36 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_35 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_35;

architecture SYN_ARCH2 of ND2_35 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_34 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_34;

architecture SYN_ARCH2 of ND2_34 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_33 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_33;

architecture SYN_ARCH2 of ND2_33 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_32 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_32;

architecture SYN_ARCH2 of ND2_32 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_31 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_31;

architecture SYN_ARCH2 of ND2_31 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_30 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_30;

architecture SYN_ARCH2 of ND2_30 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_29 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_29;

architecture SYN_ARCH2 of ND2_29 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_28 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_28;

architecture SYN_ARCH2 of ND2_28 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_27 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_27;

architecture SYN_ARCH2 of ND2_27 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_26 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_26;

architecture SYN_ARCH2 of ND2_26 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_25 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_25;

architecture SYN_ARCH2 of ND2_25 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_24 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_24;

architecture SYN_ARCH2 of ND2_24 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_23 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_23;

architecture SYN_ARCH2 of ND2_23 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_22 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_22;

architecture SYN_ARCH2 of ND2_22 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_21 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_21;

architecture SYN_ARCH2 of ND2_21 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_20 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_20;

architecture SYN_ARCH2 of ND2_20 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_19 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_19;

architecture SYN_ARCH2 of ND2_19 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_18 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_18;

architecture SYN_ARCH2 of ND2_18 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_17 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_17;

architecture SYN_ARCH2 of ND2_17 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_16 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_16;

architecture SYN_ARCH2 of ND2_16 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_15 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_15;

architecture SYN_ARCH2 of ND2_15 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_14 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_14;

architecture SYN_ARCH2 of ND2_14 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_13 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_13;

architecture SYN_ARCH2 of ND2_13 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_12 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_12;

architecture SYN_ARCH2 of ND2_12 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_11 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_11;

architecture SYN_ARCH2 of ND2_11 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_10 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_10;

architecture SYN_ARCH2 of ND2_10 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_9 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_9;

architecture SYN_ARCH2 of ND2_9 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_8 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_8;

architecture SYN_ARCH2 of ND2_8 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_7 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_7;

architecture SYN_ARCH2 of ND2_7 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_6 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_6;

architecture SYN_ARCH2 of ND2_6 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_5 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_5;

architecture SYN_ARCH2 of ND2_5 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_4 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_4;

architecture SYN_ARCH2 of ND2_4 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_3 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_3;

architecture SYN_ARCH2 of ND2_3 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_2 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_2;

architecture SYN_ARCH2 of ND2_2 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_1 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_1;

architecture SYN_ARCH2 of ND2_1 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_255 is

   port( A : in std_logic;  Y : out std_logic);

end IV_255;

architecture SYN_BEHAVIORAL of IV_255 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_254 is

   port( A : in std_logic;  Y : out std_logic);

end IV_254;

architecture SYN_BEHAVIORAL of IV_254 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_253 is

   port( A : in std_logic;  Y : out std_logic);

end IV_253;

architecture SYN_BEHAVIORAL of IV_253 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_252 is

   port( A : in std_logic;  Y : out std_logic);

end IV_252;

architecture SYN_BEHAVIORAL of IV_252 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_251 is

   port( A : in std_logic;  Y : out std_logic);

end IV_251;

architecture SYN_BEHAVIORAL of IV_251 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_250 is

   port( A : in std_logic;  Y : out std_logic);

end IV_250;

architecture SYN_BEHAVIORAL of IV_250 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_249 is

   port( A : in std_logic;  Y : out std_logic);

end IV_249;

architecture SYN_BEHAVIORAL of IV_249 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_248 is

   port( A : in std_logic;  Y : out std_logic);

end IV_248;

architecture SYN_BEHAVIORAL of IV_248 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_247 is

   port( A : in std_logic;  Y : out std_logic);

end IV_247;

architecture SYN_BEHAVIORAL of IV_247 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_246 is

   port( A : in std_logic;  Y : out std_logic);

end IV_246;

architecture SYN_BEHAVIORAL of IV_246 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_245 is

   port( A : in std_logic;  Y : out std_logic);

end IV_245;

architecture SYN_BEHAVIORAL of IV_245 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_244 is

   port( A : in std_logic;  Y : out std_logic);

end IV_244;

architecture SYN_BEHAVIORAL of IV_244 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_243 is

   port( A : in std_logic;  Y : out std_logic);

end IV_243;

architecture SYN_BEHAVIORAL of IV_243 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_242 is

   port( A : in std_logic;  Y : out std_logic);

end IV_242;

architecture SYN_BEHAVIORAL of IV_242 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_241 is

   port( A : in std_logic;  Y : out std_logic);

end IV_241;

architecture SYN_BEHAVIORAL of IV_241 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_240 is

   port( A : in std_logic;  Y : out std_logic);

end IV_240;

architecture SYN_BEHAVIORAL of IV_240 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_239 is

   port( A : in std_logic;  Y : out std_logic);

end IV_239;

architecture SYN_BEHAVIORAL of IV_239 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_238 is

   port( A : in std_logic;  Y : out std_logic);

end IV_238;

architecture SYN_BEHAVIORAL of IV_238 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_237 is

   port( A : in std_logic;  Y : out std_logic);

end IV_237;

architecture SYN_BEHAVIORAL of IV_237 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_236 is

   port( A : in std_logic;  Y : out std_logic);

end IV_236;

architecture SYN_BEHAVIORAL of IV_236 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_235 is

   port( A : in std_logic;  Y : out std_logic);

end IV_235;

architecture SYN_BEHAVIORAL of IV_235 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_234 is

   port( A : in std_logic;  Y : out std_logic);

end IV_234;

architecture SYN_BEHAVIORAL of IV_234 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_233 is

   port( A : in std_logic;  Y : out std_logic);

end IV_233;

architecture SYN_BEHAVIORAL of IV_233 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_232 is

   port( A : in std_logic;  Y : out std_logic);

end IV_232;

architecture SYN_BEHAVIORAL of IV_232 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_231 is

   port( A : in std_logic;  Y : out std_logic);

end IV_231;

architecture SYN_BEHAVIORAL of IV_231 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_230 is

   port( A : in std_logic;  Y : out std_logic);

end IV_230;

architecture SYN_BEHAVIORAL of IV_230 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_229 is

   port( A : in std_logic;  Y : out std_logic);

end IV_229;

architecture SYN_BEHAVIORAL of IV_229 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_228 is

   port( A : in std_logic;  Y : out std_logic);

end IV_228;

architecture SYN_BEHAVIORAL of IV_228 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_227 is

   port( A : in std_logic;  Y : out std_logic);

end IV_227;

architecture SYN_BEHAVIORAL of IV_227 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_226 is

   port( A : in std_logic;  Y : out std_logic);

end IV_226;

architecture SYN_BEHAVIORAL of IV_226 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_225 is

   port( A : in std_logic;  Y : out std_logic);

end IV_225;

architecture SYN_BEHAVIORAL of IV_225 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_224 is

   port( A : in std_logic;  Y : out std_logic);

end IV_224;

architecture SYN_BEHAVIORAL of IV_224 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_223 is

   port( A : in std_logic;  Y : out std_logic);

end IV_223;

architecture SYN_BEHAVIORAL of IV_223 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_222 is

   port( A : in std_logic;  Y : out std_logic);

end IV_222;

architecture SYN_BEHAVIORAL of IV_222 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_221 is

   port( A : in std_logic;  Y : out std_logic);

end IV_221;

architecture SYN_BEHAVIORAL of IV_221 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_220 is

   port( A : in std_logic;  Y : out std_logic);

end IV_220;

architecture SYN_BEHAVIORAL of IV_220 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_219 is

   port( A : in std_logic;  Y : out std_logic);

end IV_219;

architecture SYN_BEHAVIORAL of IV_219 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_218 is

   port( A : in std_logic;  Y : out std_logic);

end IV_218;

architecture SYN_BEHAVIORAL of IV_218 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_217 is

   port( A : in std_logic;  Y : out std_logic);

end IV_217;

architecture SYN_BEHAVIORAL of IV_217 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_216 is

   port( A : in std_logic;  Y : out std_logic);

end IV_216;

architecture SYN_BEHAVIORAL of IV_216 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_215 is

   port( A : in std_logic;  Y : out std_logic);

end IV_215;

architecture SYN_BEHAVIORAL of IV_215 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_214 is

   port( A : in std_logic;  Y : out std_logic);

end IV_214;

architecture SYN_BEHAVIORAL of IV_214 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_213 is

   port( A : in std_logic;  Y : out std_logic);

end IV_213;

architecture SYN_BEHAVIORAL of IV_213 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_212 is

   port( A : in std_logic;  Y : out std_logic);

end IV_212;

architecture SYN_BEHAVIORAL of IV_212 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_211 is

   port( A : in std_logic;  Y : out std_logic);

end IV_211;

architecture SYN_BEHAVIORAL of IV_211 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_210 is

   port( A : in std_logic;  Y : out std_logic);

end IV_210;

architecture SYN_BEHAVIORAL of IV_210 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_209 is

   port( A : in std_logic;  Y : out std_logic);

end IV_209;

architecture SYN_BEHAVIORAL of IV_209 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_208 is

   port( A : in std_logic;  Y : out std_logic);

end IV_208;

architecture SYN_BEHAVIORAL of IV_208 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_207 is

   port( A : in std_logic;  Y : out std_logic);

end IV_207;

architecture SYN_BEHAVIORAL of IV_207 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_206 is

   port( A : in std_logic;  Y : out std_logic);

end IV_206;

architecture SYN_BEHAVIORAL of IV_206 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_205 is

   port( A : in std_logic;  Y : out std_logic);

end IV_205;

architecture SYN_BEHAVIORAL of IV_205 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_204 is

   port( A : in std_logic;  Y : out std_logic);

end IV_204;

architecture SYN_BEHAVIORAL of IV_204 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_203 is

   port( A : in std_logic;  Y : out std_logic);

end IV_203;

architecture SYN_BEHAVIORAL of IV_203 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_202 is

   port( A : in std_logic;  Y : out std_logic);

end IV_202;

architecture SYN_BEHAVIORAL of IV_202 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_201 is

   port( A : in std_logic;  Y : out std_logic);

end IV_201;

architecture SYN_BEHAVIORAL of IV_201 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_200 is

   port( A : in std_logic;  Y : out std_logic);

end IV_200;

architecture SYN_BEHAVIORAL of IV_200 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_199 is

   port( A : in std_logic;  Y : out std_logic);

end IV_199;

architecture SYN_BEHAVIORAL of IV_199 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_198 is

   port( A : in std_logic;  Y : out std_logic);

end IV_198;

architecture SYN_BEHAVIORAL of IV_198 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_197 is

   port( A : in std_logic;  Y : out std_logic);

end IV_197;

architecture SYN_BEHAVIORAL of IV_197 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_196 is

   port( A : in std_logic;  Y : out std_logic);

end IV_196;

architecture SYN_BEHAVIORAL of IV_196 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_195 is

   port( A : in std_logic;  Y : out std_logic);

end IV_195;

architecture SYN_BEHAVIORAL of IV_195 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_194 is

   port( A : in std_logic;  Y : out std_logic);

end IV_194;

architecture SYN_BEHAVIORAL of IV_194 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_193 is

   port( A : in std_logic;  Y : out std_logic);

end IV_193;

architecture SYN_BEHAVIORAL of IV_193 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_192 is

   port( A : in std_logic;  Y : out std_logic);

end IV_192;

architecture SYN_BEHAVIORAL of IV_192 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_191 is

   port( A : in std_logic;  Y : out std_logic);

end IV_191;

architecture SYN_BEHAVIORAL of IV_191 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_190 is

   port( A : in std_logic;  Y : out std_logic);

end IV_190;

architecture SYN_BEHAVIORAL of IV_190 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_189 is

   port( A : in std_logic;  Y : out std_logic);

end IV_189;

architecture SYN_BEHAVIORAL of IV_189 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_188 is

   port( A : in std_logic;  Y : out std_logic);

end IV_188;

architecture SYN_BEHAVIORAL of IV_188 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_187 is

   port( A : in std_logic;  Y : out std_logic);

end IV_187;

architecture SYN_BEHAVIORAL of IV_187 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_186 is

   port( A : in std_logic;  Y : out std_logic);

end IV_186;

architecture SYN_BEHAVIORAL of IV_186 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_185 is

   port( A : in std_logic;  Y : out std_logic);

end IV_185;

architecture SYN_BEHAVIORAL of IV_185 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_184 is

   port( A : in std_logic;  Y : out std_logic);

end IV_184;

architecture SYN_BEHAVIORAL of IV_184 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_183 is

   port( A : in std_logic;  Y : out std_logic);

end IV_183;

architecture SYN_BEHAVIORAL of IV_183 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_182 is

   port( A : in std_logic;  Y : out std_logic);

end IV_182;

architecture SYN_BEHAVIORAL of IV_182 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_181 is

   port( A : in std_logic;  Y : out std_logic);

end IV_181;

architecture SYN_BEHAVIORAL of IV_181 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_180 is

   port( A : in std_logic;  Y : out std_logic);

end IV_180;

architecture SYN_BEHAVIORAL of IV_180 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_179 is

   port( A : in std_logic;  Y : out std_logic);

end IV_179;

architecture SYN_BEHAVIORAL of IV_179 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_178 is

   port( A : in std_logic;  Y : out std_logic);

end IV_178;

architecture SYN_BEHAVIORAL of IV_178 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_177 is

   port( A : in std_logic;  Y : out std_logic);

end IV_177;

architecture SYN_BEHAVIORAL of IV_177 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_176 is

   port( A : in std_logic;  Y : out std_logic);

end IV_176;

architecture SYN_BEHAVIORAL of IV_176 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_175 is

   port( A : in std_logic;  Y : out std_logic);

end IV_175;

architecture SYN_BEHAVIORAL of IV_175 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_174 is

   port( A : in std_logic;  Y : out std_logic);

end IV_174;

architecture SYN_BEHAVIORAL of IV_174 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_173 is

   port( A : in std_logic;  Y : out std_logic);

end IV_173;

architecture SYN_BEHAVIORAL of IV_173 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_172 is

   port( A : in std_logic;  Y : out std_logic);

end IV_172;

architecture SYN_BEHAVIORAL of IV_172 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_171 is

   port( A : in std_logic;  Y : out std_logic);

end IV_171;

architecture SYN_BEHAVIORAL of IV_171 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_170 is

   port( A : in std_logic;  Y : out std_logic);

end IV_170;

architecture SYN_BEHAVIORAL of IV_170 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_169 is

   port( A : in std_logic;  Y : out std_logic);

end IV_169;

architecture SYN_BEHAVIORAL of IV_169 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_168 is

   port( A : in std_logic;  Y : out std_logic);

end IV_168;

architecture SYN_BEHAVIORAL of IV_168 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_167 is

   port( A : in std_logic;  Y : out std_logic);

end IV_167;

architecture SYN_BEHAVIORAL of IV_167 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_166 is

   port( A : in std_logic;  Y : out std_logic);

end IV_166;

architecture SYN_BEHAVIORAL of IV_166 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_165 is

   port( A : in std_logic;  Y : out std_logic);

end IV_165;

architecture SYN_BEHAVIORAL of IV_165 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_164 is

   port( A : in std_logic;  Y : out std_logic);

end IV_164;

architecture SYN_BEHAVIORAL of IV_164 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_163 is

   port( A : in std_logic;  Y : out std_logic);

end IV_163;

architecture SYN_BEHAVIORAL of IV_163 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_162 is

   port( A : in std_logic;  Y : out std_logic);

end IV_162;

architecture SYN_BEHAVIORAL of IV_162 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_161 is

   port( A : in std_logic;  Y : out std_logic);

end IV_161;

architecture SYN_BEHAVIORAL of IV_161 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_160 is

   port( A : in std_logic;  Y : out std_logic);

end IV_160;

architecture SYN_BEHAVIORAL of IV_160 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_159 is

   port( A : in std_logic;  Y : out std_logic);

end IV_159;

architecture SYN_BEHAVIORAL of IV_159 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_158 is

   port( A : in std_logic;  Y : out std_logic);

end IV_158;

architecture SYN_BEHAVIORAL of IV_158 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_157 is

   port( A : in std_logic;  Y : out std_logic);

end IV_157;

architecture SYN_BEHAVIORAL of IV_157 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_156 is

   port( A : in std_logic;  Y : out std_logic);

end IV_156;

architecture SYN_BEHAVIORAL of IV_156 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_155 is

   port( A : in std_logic;  Y : out std_logic);

end IV_155;

architecture SYN_BEHAVIORAL of IV_155 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_154 is

   port( A : in std_logic;  Y : out std_logic);

end IV_154;

architecture SYN_BEHAVIORAL of IV_154 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_153 is

   port( A : in std_logic;  Y : out std_logic);

end IV_153;

architecture SYN_BEHAVIORAL of IV_153 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_152 is

   port( A : in std_logic;  Y : out std_logic);

end IV_152;

architecture SYN_BEHAVIORAL of IV_152 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_151 is

   port( A : in std_logic;  Y : out std_logic);

end IV_151;

architecture SYN_BEHAVIORAL of IV_151 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_150 is

   port( A : in std_logic;  Y : out std_logic);

end IV_150;

architecture SYN_BEHAVIORAL of IV_150 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_149 is

   port( A : in std_logic;  Y : out std_logic);

end IV_149;

architecture SYN_BEHAVIORAL of IV_149 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_148 is

   port( A : in std_logic;  Y : out std_logic);

end IV_148;

architecture SYN_BEHAVIORAL of IV_148 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_147 is

   port( A : in std_logic;  Y : out std_logic);

end IV_147;

architecture SYN_BEHAVIORAL of IV_147 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_146 is

   port( A : in std_logic;  Y : out std_logic);

end IV_146;

architecture SYN_BEHAVIORAL of IV_146 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_145 is

   port( A : in std_logic;  Y : out std_logic);

end IV_145;

architecture SYN_BEHAVIORAL of IV_145 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_144 is

   port( A : in std_logic;  Y : out std_logic);

end IV_144;

architecture SYN_BEHAVIORAL of IV_144 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_143 is

   port( A : in std_logic;  Y : out std_logic);

end IV_143;

architecture SYN_BEHAVIORAL of IV_143 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_142 is

   port( A : in std_logic;  Y : out std_logic);

end IV_142;

architecture SYN_BEHAVIORAL of IV_142 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_141 is

   port( A : in std_logic;  Y : out std_logic);

end IV_141;

architecture SYN_BEHAVIORAL of IV_141 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_140 is

   port( A : in std_logic;  Y : out std_logic);

end IV_140;

architecture SYN_BEHAVIORAL of IV_140 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_139 is

   port( A : in std_logic;  Y : out std_logic);

end IV_139;

architecture SYN_BEHAVIORAL of IV_139 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_138 is

   port( A : in std_logic;  Y : out std_logic);

end IV_138;

architecture SYN_BEHAVIORAL of IV_138 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_137 is

   port( A : in std_logic;  Y : out std_logic);

end IV_137;

architecture SYN_BEHAVIORAL of IV_137 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_136 is

   port( A : in std_logic;  Y : out std_logic);

end IV_136;

architecture SYN_BEHAVIORAL of IV_136 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_135 is

   port( A : in std_logic;  Y : out std_logic);

end IV_135;

architecture SYN_BEHAVIORAL of IV_135 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_134 is

   port( A : in std_logic;  Y : out std_logic);

end IV_134;

architecture SYN_BEHAVIORAL of IV_134 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_133 is

   port( A : in std_logic;  Y : out std_logic);

end IV_133;

architecture SYN_BEHAVIORAL of IV_133 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_132 is

   port( A : in std_logic;  Y : out std_logic);

end IV_132;

architecture SYN_BEHAVIORAL of IV_132 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_131 is

   port( A : in std_logic;  Y : out std_logic);

end IV_131;

architecture SYN_BEHAVIORAL of IV_131 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_130 is

   port( A : in std_logic;  Y : out std_logic);

end IV_130;

architecture SYN_BEHAVIORAL of IV_130 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_129 is

   port( A : in std_logic;  Y : out std_logic);

end IV_129;

architecture SYN_BEHAVIORAL of IV_129 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_128 is

   port( A : in std_logic;  Y : out std_logic);

end IV_128;

architecture SYN_BEHAVIORAL of IV_128 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_127 is

   port( A : in std_logic;  Y : out std_logic);

end IV_127;

architecture SYN_BEHAVIORAL of IV_127 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_126 is

   port( A : in std_logic;  Y : out std_logic);

end IV_126;

architecture SYN_BEHAVIORAL of IV_126 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_125 is

   port( A : in std_logic;  Y : out std_logic);

end IV_125;

architecture SYN_BEHAVIORAL of IV_125 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_124 is

   port( A : in std_logic;  Y : out std_logic);

end IV_124;

architecture SYN_BEHAVIORAL of IV_124 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_123 is

   port( A : in std_logic;  Y : out std_logic);

end IV_123;

architecture SYN_BEHAVIORAL of IV_123 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_122 is

   port( A : in std_logic;  Y : out std_logic);

end IV_122;

architecture SYN_BEHAVIORAL of IV_122 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_121 is

   port( A : in std_logic;  Y : out std_logic);

end IV_121;

architecture SYN_BEHAVIORAL of IV_121 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_120 is

   port( A : in std_logic;  Y : out std_logic);

end IV_120;

architecture SYN_BEHAVIORAL of IV_120 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_119 is

   port( A : in std_logic;  Y : out std_logic);

end IV_119;

architecture SYN_BEHAVIORAL of IV_119 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_118 is

   port( A : in std_logic;  Y : out std_logic);

end IV_118;

architecture SYN_BEHAVIORAL of IV_118 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_117 is

   port( A : in std_logic;  Y : out std_logic);

end IV_117;

architecture SYN_BEHAVIORAL of IV_117 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_116 is

   port( A : in std_logic;  Y : out std_logic);

end IV_116;

architecture SYN_BEHAVIORAL of IV_116 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_115 is

   port( A : in std_logic;  Y : out std_logic);

end IV_115;

architecture SYN_BEHAVIORAL of IV_115 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_114 is

   port( A : in std_logic;  Y : out std_logic);

end IV_114;

architecture SYN_BEHAVIORAL of IV_114 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_113 is

   port( A : in std_logic;  Y : out std_logic);

end IV_113;

architecture SYN_BEHAVIORAL of IV_113 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_112 is

   port( A : in std_logic;  Y : out std_logic);

end IV_112;

architecture SYN_BEHAVIORAL of IV_112 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_111 is

   port( A : in std_logic;  Y : out std_logic);

end IV_111;

architecture SYN_BEHAVIORAL of IV_111 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_110 is

   port( A : in std_logic;  Y : out std_logic);

end IV_110;

architecture SYN_BEHAVIORAL of IV_110 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_109 is

   port( A : in std_logic;  Y : out std_logic);

end IV_109;

architecture SYN_BEHAVIORAL of IV_109 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_108 is

   port( A : in std_logic;  Y : out std_logic);

end IV_108;

architecture SYN_BEHAVIORAL of IV_108 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_107 is

   port( A : in std_logic;  Y : out std_logic);

end IV_107;

architecture SYN_BEHAVIORAL of IV_107 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_106 is

   port( A : in std_logic;  Y : out std_logic);

end IV_106;

architecture SYN_BEHAVIORAL of IV_106 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_105 is

   port( A : in std_logic;  Y : out std_logic);

end IV_105;

architecture SYN_BEHAVIORAL of IV_105 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_104 is

   port( A : in std_logic;  Y : out std_logic);

end IV_104;

architecture SYN_BEHAVIORAL of IV_104 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_103 is

   port( A : in std_logic;  Y : out std_logic);

end IV_103;

architecture SYN_BEHAVIORAL of IV_103 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_102 is

   port( A : in std_logic;  Y : out std_logic);

end IV_102;

architecture SYN_BEHAVIORAL of IV_102 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_101 is

   port( A : in std_logic;  Y : out std_logic);

end IV_101;

architecture SYN_BEHAVIORAL of IV_101 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_100 is

   port( A : in std_logic;  Y : out std_logic);

end IV_100;

architecture SYN_BEHAVIORAL of IV_100 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_99 is

   port( A : in std_logic;  Y : out std_logic);

end IV_99;

architecture SYN_BEHAVIORAL of IV_99 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_98 is

   port( A : in std_logic;  Y : out std_logic);

end IV_98;

architecture SYN_BEHAVIORAL of IV_98 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_97 is

   port( A : in std_logic;  Y : out std_logic);

end IV_97;

architecture SYN_BEHAVIORAL of IV_97 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_96 is

   port( A : in std_logic;  Y : out std_logic);

end IV_96;

architecture SYN_BEHAVIORAL of IV_96 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_95 is

   port( A : in std_logic;  Y : out std_logic);

end IV_95;

architecture SYN_BEHAVIORAL of IV_95 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_94 is

   port( A : in std_logic;  Y : out std_logic);

end IV_94;

architecture SYN_BEHAVIORAL of IV_94 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_93 is

   port( A : in std_logic;  Y : out std_logic);

end IV_93;

architecture SYN_BEHAVIORAL of IV_93 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_92 is

   port( A : in std_logic;  Y : out std_logic);

end IV_92;

architecture SYN_BEHAVIORAL of IV_92 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_91 is

   port( A : in std_logic;  Y : out std_logic);

end IV_91;

architecture SYN_BEHAVIORAL of IV_91 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_90 is

   port( A : in std_logic;  Y : out std_logic);

end IV_90;

architecture SYN_BEHAVIORAL of IV_90 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_89 is

   port( A : in std_logic;  Y : out std_logic);

end IV_89;

architecture SYN_BEHAVIORAL of IV_89 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_88 is

   port( A : in std_logic;  Y : out std_logic);

end IV_88;

architecture SYN_BEHAVIORAL of IV_88 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_87 is

   port( A : in std_logic;  Y : out std_logic);

end IV_87;

architecture SYN_BEHAVIORAL of IV_87 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_86 is

   port( A : in std_logic;  Y : out std_logic);

end IV_86;

architecture SYN_BEHAVIORAL of IV_86 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_85 is

   port( A : in std_logic;  Y : out std_logic);

end IV_85;

architecture SYN_BEHAVIORAL of IV_85 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_84 is

   port( A : in std_logic;  Y : out std_logic);

end IV_84;

architecture SYN_BEHAVIORAL of IV_84 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_83 is

   port( A : in std_logic;  Y : out std_logic);

end IV_83;

architecture SYN_BEHAVIORAL of IV_83 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_82 is

   port( A : in std_logic;  Y : out std_logic);

end IV_82;

architecture SYN_BEHAVIORAL of IV_82 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_81 is

   port( A : in std_logic;  Y : out std_logic);

end IV_81;

architecture SYN_BEHAVIORAL of IV_81 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_80 is

   port( A : in std_logic;  Y : out std_logic);

end IV_80;

architecture SYN_BEHAVIORAL of IV_80 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_79 is

   port( A : in std_logic;  Y : out std_logic);

end IV_79;

architecture SYN_BEHAVIORAL of IV_79 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_78 is

   port( A : in std_logic;  Y : out std_logic);

end IV_78;

architecture SYN_BEHAVIORAL of IV_78 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_77 is

   port( A : in std_logic;  Y : out std_logic);

end IV_77;

architecture SYN_BEHAVIORAL of IV_77 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_76 is

   port( A : in std_logic;  Y : out std_logic);

end IV_76;

architecture SYN_BEHAVIORAL of IV_76 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_75 is

   port( A : in std_logic;  Y : out std_logic);

end IV_75;

architecture SYN_BEHAVIORAL of IV_75 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_74 is

   port( A : in std_logic;  Y : out std_logic);

end IV_74;

architecture SYN_BEHAVIORAL of IV_74 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_73 is

   port( A : in std_logic;  Y : out std_logic);

end IV_73;

architecture SYN_BEHAVIORAL of IV_73 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_72 is

   port( A : in std_logic;  Y : out std_logic);

end IV_72;

architecture SYN_BEHAVIORAL of IV_72 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_71 is

   port( A : in std_logic;  Y : out std_logic);

end IV_71;

architecture SYN_BEHAVIORAL of IV_71 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_70 is

   port( A : in std_logic;  Y : out std_logic);

end IV_70;

architecture SYN_BEHAVIORAL of IV_70 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_69 is

   port( A : in std_logic;  Y : out std_logic);

end IV_69;

architecture SYN_BEHAVIORAL of IV_69 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_68 is

   port( A : in std_logic;  Y : out std_logic);

end IV_68;

architecture SYN_BEHAVIORAL of IV_68 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_67 is

   port( A : in std_logic;  Y : out std_logic);

end IV_67;

architecture SYN_BEHAVIORAL of IV_67 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_66 is

   port( A : in std_logic;  Y : out std_logic);

end IV_66;

architecture SYN_BEHAVIORAL of IV_66 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_65 is

   port( A : in std_logic;  Y : out std_logic);

end IV_65;

architecture SYN_BEHAVIORAL of IV_65 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_64 is

   port( A : in std_logic;  Y : out std_logic);

end IV_64;

architecture SYN_BEHAVIORAL of IV_64 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_63 is

   port( A : in std_logic;  Y : out std_logic);

end IV_63;

architecture SYN_BEHAVIORAL of IV_63 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_62 is

   port( A : in std_logic;  Y : out std_logic);

end IV_62;

architecture SYN_BEHAVIORAL of IV_62 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_61 is

   port( A : in std_logic;  Y : out std_logic);

end IV_61;

architecture SYN_BEHAVIORAL of IV_61 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_60 is

   port( A : in std_logic;  Y : out std_logic);

end IV_60;

architecture SYN_BEHAVIORAL of IV_60 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_59 is

   port( A : in std_logic;  Y : out std_logic);

end IV_59;

architecture SYN_BEHAVIORAL of IV_59 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_58 is

   port( A : in std_logic;  Y : out std_logic);

end IV_58;

architecture SYN_BEHAVIORAL of IV_58 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_57 is

   port( A : in std_logic;  Y : out std_logic);

end IV_57;

architecture SYN_BEHAVIORAL of IV_57 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_56 is

   port( A : in std_logic;  Y : out std_logic);

end IV_56;

architecture SYN_BEHAVIORAL of IV_56 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_55 is

   port( A : in std_logic;  Y : out std_logic);

end IV_55;

architecture SYN_BEHAVIORAL of IV_55 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_54 is

   port( A : in std_logic;  Y : out std_logic);

end IV_54;

architecture SYN_BEHAVIORAL of IV_54 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_53 is

   port( A : in std_logic;  Y : out std_logic);

end IV_53;

architecture SYN_BEHAVIORAL of IV_53 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_52 is

   port( A : in std_logic;  Y : out std_logic);

end IV_52;

architecture SYN_BEHAVIORAL of IV_52 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_51 is

   port( A : in std_logic;  Y : out std_logic);

end IV_51;

architecture SYN_BEHAVIORAL of IV_51 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_50 is

   port( A : in std_logic;  Y : out std_logic);

end IV_50;

architecture SYN_BEHAVIORAL of IV_50 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_49 is

   port( A : in std_logic;  Y : out std_logic);

end IV_49;

architecture SYN_BEHAVIORAL of IV_49 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_48 is

   port( A : in std_logic;  Y : out std_logic);

end IV_48;

architecture SYN_BEHAVIORAL of IV_48 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_47 is

   port( A : in std_logic;  Y : out std_logic);

end IV_47;

architecture SYN_BEHAVIORAL of IV_47 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_46 is

   port( A : in std_logic;  Y : out std_logic);

end IV_46;

architecture SYN_BEHAVIORAL of IV_46 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_45 is

   port( A : in std_logic;  Y : out std_logic);

end IV_45;

architecture SYN_BEHAVIORAL of IV_45 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_44 is

   port( A : in std_logic;  Y : out std_logic);

end IV_44;

architecture SYN_BEHAVIORAL of IV_44 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_43 is

   port( A : in std_logic;  Y : out std_logic);

end IV_43;

architecture SYN_BEHAVIORAL of IV_43 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_42 is

   port( A : in std_logic;  Y : out std_logic);

end IV_42;

architecture SYN_BEHAVIORAL of IV_42 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_41 is

   port( A : in std_logic;  Y : out std_logic);

end IV_41;

architecture SYN_BEHAVIORAL of IV_41 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_40 is

   port( A : in std_logic;  Y : out std_logic);

end IV_40;

architecture SYN_BEHAVIORAL of IV_40 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_39 is

   port( A : in std_logic;  Y : out std_logic);

end IV_39;

architecture SYN_BEHAVIORAL of IV_39 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_38 is

   port( A : in std_logic;  Y : out std_logic);

end IV_38;

architecture SYN_BEHAVIORAL of IV_38 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_37 is

   port( A : in std_logic;  Y : out std_logic);

end IV_37;

architecture SYN_BEHAVIORAL of IV_37 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_36 is

   port( A : in std_logic;  Y : out std_logic);

end IV_36;

architecture SYN_BEHAVIORAL of IV_36 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_35 is

   port( A : in std_logic;  Y : out std_logic);

end IV_35;

architecture SYN_BEHAVIORAL of IV_35 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_34 is

   port( A : in std_logic;  Y : out std_logic);

end IV_34;

architecture SYN_BEHAVIORAL of IV_34 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_33 is

   port( A : in std_logic;  Y : out std_logic);

end IV_33;

architecture SYN_BEHAVIORAL of IV_33 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_32 is

   port( A : in std_logic;  Y : out std_logic);

end IV_32;

architecture SYN_BEHAVIORAL of IV_32 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_31 is

   port( A : in std_logic;  Y : out std_logic);

end IV_31;

architecture SYN_BEHAVIORAL of IV_31 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_30 is

   port( A : in std_logic;  Y : out std_logic);

end IV_30;

architecture SYN_BEHAVIORAL of IV_30 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_29 is

   port( A : in std_logic;  Y : out std_logic);

end IV_29;

architecture SYN_BEHAVIORAL of IV_29 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_28 is

   port( A : in std_logic;  Y : out std_logic);

end IV_28;

architecture SYN_BEHAVIORAL of IV_28 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_27 is

   port( A : in std_logic;  Y : out std_logic);

end IV_27;

architecture SYN_BEHAVIORAL of IV_27 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_26 is

   port( A : in std_logic;  Y : out std_logic);

end IV_26;

architecture SYN_BEHAVIORAL of IV_26 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_25 is

   port( A : in std_logic;  Y : out std_logic);

end IV_25;

architecture SYN_BEHAVIORAL of IV_25 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_24 is

   port( A : in std_logic;  Y : out std_logic);

end IV_24;

architecture SYN_BEHAVIORAL of IV_24 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_23 is

   port( A : in std_logic;  Y : out std_logic);

end IV_23;

architecture SYN_BEHAVIORAL of IV_23 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_22 is

   port( A : in std_logic;  Y : out std_logic);

end IV_22;

architecture SYN_BEHAVIORAL of IV_22 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_21 is

   port( A : in std_logic;  Y : out std_logic);

end IV_21;

architecture SYN_BEHAVIORAL of IV_21 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_20 is

   port( A : in std_logic;  Y : out std_logic);

end IV_20;

architecture SYN_BEHAVIORAL of IV_20 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_19 is

   port( A : in std_logic;  Y : out std_logic);

end IV_19;

architecture SYN_BEHAVIORAL of IV_19 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_18 is

   port( A : in std_logic;  Y : out std_logic);

end IV_18;

architecture SYN_BEHAVIORAL of IV_18 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_17 is

   port( A : in std_logic;  Y : out std_logic);

end IV_17;

architecture SYN_BEHAVIORAL of IV_17 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_16 is

   port( A : in std_logic;  Y : out std_logic);

end IV_16;

architecture SYN_BEHAVIORAL of IV_16 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_15 is

   port( A : in std_logic;  Y : out std_logic);

end IV_15;

architecture SYN_BEHAVIORAL of IV_15 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_14 is

   port( A : in std_logic;  Y : out std_logic);

end IV_14;

architecture SYN_BEHAVIORAL of IV_14 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_13 is

   port( A : in std_logic;  Y : out std_logic);

end IV_13;

architecture SYN_BEHAVIORAL of IV_13 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_12 is

   port( A : in std_logic;  Y : out std_logic);

end IV_12;

architecture SYN_BEHAVIORAL of IV_12 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_11 is

   port( A : in std_logic;  Y : out std_logic);

end IV_11;

architecture SYN_BEHAVIORAL of IV_11 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_10 is

   port( A : in std_logic;  Y : out std_logic);

end IV_10;

architecture SYN_BEHAVIORAL of IV_10 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_9 is

   port( A : in std_logic;  Y : out std_logic);

end IV_9;

architecture SYN_BEHAVIORAL of IV_9 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_8 is

   port( A : in std_logic;  Y : out std_logic);

end IV_8;

architecture SYN_BEHAVIORAL of IV_8 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_7 is

   port( A : in std_logic;  Y : out std_logic);

end IV_7;

architecture SYN_BEHAVIORAL of IV_7 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_6 is

   port( A : in std_logic;  Y : out std_logic);

end IV_6;

architecture SYN_BEHAVIORAL of IV_6 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_5 is

   port( A : in std_logic;  Y : out std_logic);

end IV_5;

architecture SYN_BEHAVIORAL of IV_5 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_4 is

   port( A : in std_logic;  Y : out std_logic);

end IV_4;

architecture SYN_BEHAVIORAL of IV_4 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_3 is

   port( A : in std_logic;  Y : out std_logic);

end IV_3;

architecture SYN_BEHAVIORAL of IV_3 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_2 is

   port( A : in std_logic;  Y : out std_logic);

end IV_2;

architecture SYN_BEHAVIORAL of IV_2 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_1 is

   port( A : in std_logic;  Y : out std_logic);

end IV_1;

architecture SYN_BEHAVIORAL of IV_1 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_255 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_255;

architecture SYN_STRUCTURAL of MUX21_255 is

   component ND2_763
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_764
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_765
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_255
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_255 port map( A => S, Y => SB);
   UND1 : ND2_765 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_764 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_763 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_254 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_254;

architecture SYN_STRUCTURAL of MUX21_254 is

   component ND2_760
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_761
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_762
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_254
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_254 port map( A => S, Y => SB);
   UND1 : ND2_762 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_761 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_760 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_253 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_253;

architecture SYN_STRUCTURAL of MUX21_253 is

   component ND2_757
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_758
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_759
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_253
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_253 port map( A => S, Y => SB);
   UND1 : ND2_759 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_758 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_757 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_252 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_252;

architecture SYN_STRUCTURAL of MUX21_252 is

   component ND2_754
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_755
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_756
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_252
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_252 port map( A => S, Y => SB);
   UND1 : ND2_756 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_755 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_754 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_251 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_251;

architecture SYN_STRUCTURAL of MUX21_251 is

   component ND2_751
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_752
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_753
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_251
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_251 port map( A => S, Y => SB);
   UND1 : ND2_753 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_752 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_751 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_250 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_250;

architecture SYN_STRUCTURAL of MUX21_250 is

   component ND2_748
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_749
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_750
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_250
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_250 port map( A => S, Y => SB);
   UND1 : ND2_750 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_749 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_748 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_249 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_249;

architecture SYN_STRUCTURAL of MUX21_249 is

   component ND2_745
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_746
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_747
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_249
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_249 port map( A => S, Y => SB);
   UND1 : ND2_747 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_746 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_745 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_248 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_248;

architecture SYN_STRUCTURAL of MUX21_248 is

   component ND2_742
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_743
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_744
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_248
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_248 port map( A => S, Y => SB);
   UND1 : ND2_744 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_743 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_742 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_247 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_247;

architecture SYN_STRUCTURAL of MUX21_247 is

   component ND2_739
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_740
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_741
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_247
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_247 port map( A => S, Y => SB);
   UND1 : ND2_741 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_740 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_739 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_246 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_246;

architecture SYN_STRUCTURAL of MUX21_246 is

   component ND2_736
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_737
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_738
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_246
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_246 port map( A => S, Y => SB);
   UND1 : ND2_738 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_737 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_736 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_245 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_245;

architecture SYN_STRUCTURAL of MUX21_245 is

   component ND2_733
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_734
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_735
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_245
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_245 port map( A => S, Y => SB);
   UND1 : ND2_735 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_734 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_733 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_244 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_244;

architecture SYN_STRUCTURAL of MUX21_244 is

   component ND2_730
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_731
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_732
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_244
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_244 port map( A => S, Y => SB);
   UND1 : ND2_732 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_731 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_730 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_243 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_243;

architecture SYN_STRUCTURAL of MUX21_243 is

   component ND2_727
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_728
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_729
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_243
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_243 port map( A => S, Y => SB);
   UND1 : ND2_729 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_728 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_727 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_242 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_242;

architecture SYN_STRUCTURAL of MUX21_242 is

   component ND2_724
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_725
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_726
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_242
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_242 port map( A => S, Y => SB);
   UND1 : ND2_726 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_725 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_724 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_241 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_241;

architecture SYN_STRUCTURAL of MUX21_241 is

   component ND2_721
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_722
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_723
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_241
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_241 port map( A => S, Y => SB);
   UND1 : ND2_723 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_722 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_721 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_240 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_240;

architecture SYN_STRUCTURAL of MUX21_240 is

   component ND2_718
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_719
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_720
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_240
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_240 port map( A => S, Y => SB);
   UND1 : ND2_720 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_719 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_718 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_239 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_239;

architecture SYN_STRUCTURAL of MUX21_239 is

   component ND2_715
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_716
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_717
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_239
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_239 port map( A => S, Y => SB);
   UND1 : ND2_717 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_716 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_715 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_238 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_238;

architecture SYN_STRUCTURAL of MUX21_238 is

   component ND2_712
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_713
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_714
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_238
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_238 port map( A => S, Y => SB);
   UND1 : ND2_714 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_713 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_712 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_237 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_237;

architecture SYN_STRUCTURAL of MUX21_237 is

   component ND2_709
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_710
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_711
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_237
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_237 port map( A => S, Y => SB);
   UND1 : ND2_711 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_710 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_709 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_236 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_236;

architecture SYN_STRUCTURAL of MUX21_236 is

   component ND2_706
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_707
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_708
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_236
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_236 port map( A => S, Y => SB);
   UND1 : ND2_708 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_707 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_706 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_235 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_235;

architecture SYN_STRUCTURAL of MUX21_235 is

   component ND2_703
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_704
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_705
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_235
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_235 port map( A => S, Y => SB);
   UND1 : ND2_705 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_704 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_703 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_234 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_234;

architecture SYN_STRUCTURAL of MUX21_234 is

   component ND2_700
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_701
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_702
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_234
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_234 port map( A => S, Y => SB);
   UND1 : ND2_702 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_701 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_700 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_233 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_233;

architecture SYN_STRUCTURAL of MUX21_233 is

   component ND2_697
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_698
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_699
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_233
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_233 port map( A => S, Y => SB);
   UND1 : ND2_699 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_698 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_697 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_232 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_232;

architecture SYN_STRUCTURAL of MUX21_232 is

   component ND2_694
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_695
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_696
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_232
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_232 port map( A => S, Y => SB);
   UND1 : ND2_696 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_695 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_694 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_231 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_231;

architecture SYN_STRUCTURAL of MUX21_231 is

   component ND2_691
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_692
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_693
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_231
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_231 port map( A => S, Y => SB);
   UND1 : ND2_693 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_692 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_691 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_230 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_230;

architecture SYN_STRUCTURAL of MUX21_230 is

   component ND2_688
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_689
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_690
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_230
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_230 port map( A => S, Y => SB);
   UND1 : ND2_690 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_689 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_688 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_229 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_229;

architecture SYN_STRUCTURAL of MUX21_229 is

   component ND2_685
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_686
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_687
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_229
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_229 port map( A => S, Y => SB);
   UND1 : ND2_687 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_686 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_685 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_228 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_228;

architecture SYN_STRUCTURAL of MUX21_228 is

   component ND2_682
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_683
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_684
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_228
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_228 port map( A => S, Y => SB);
   UND1 : ND2_684 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_683 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_682 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_227 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_227;

architecture SYN_STRUCTURAL of MUX21_227 is

   component ND2_679
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_680
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_681
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_227
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_227 port map( A => S, Y => SB);
   UND1 : ND2_681 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_680 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_679 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_226 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_226;

architecture SYN_STRUCTURAL of MUX21_226 is

   component ND2_676
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_677
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_678
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_226
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_226 port map( A => S, Y => SB);
   UND1 : ND2_678 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_677 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_676 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_225 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_225;

architecture SYN_STRUCTURAL of MUX21_225 is

   component ND2_673
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_674
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_675
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_225
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_225 port map( A => S, Y => SB);
   UND1 : ND2_675 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_674 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_673 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_224 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_224;

architecture SYN_STRUCTURAL of MUX21_224 is

   component ND2_670
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_671
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_672
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_224
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_224 port map( A => S, Y => SB);
   UND1 : ND2_672 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_671 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_670 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_223 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_223;

architecture SYN_STRUCTURAL of MUX21_223 is

   component ND2_667
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_668
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_669
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_223
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_223 port map( A => S, Y => SB);
   UND1 : ND2_669 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_668 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_667 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_222 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_222;

architecture SYN_STRUCTURAL of MUX21_222 is

   component ND2_664
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_665
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_666
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_222
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_222 port map( A => S, Y => SB);
   UND1 : ND2_666 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_665 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_664 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_221 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_221;

architecture SYN_STRUCTURAL of MUX21_221 is

   component ND2_661
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_662
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_663
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_221
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_221 port map( A => S, Y => SB);
   UND1 : ND2_663 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_662 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_661 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_220 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_220;

architecture SYN_STRUCTURAL of MUX21_220 is

   component ND2_658
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_659
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_660
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_220
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_220 port map( A => S, Y => SB);
   UND1 : ND2_660 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_659 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_658 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_219 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_219;

architecture SYN_STRUCTURAL of MUX21_219 is

   component ND2_655
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_656
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_657
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_219
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_219 port map( A => S, Y => SB);
   UND1 : ND2_657 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_656 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_655 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_218 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_218;

architecture SYN_STRUCTURAL of MUX21_218 is

   component ND2_652
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_653
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_654
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_218
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_218 port map( A => S, Y => SB);
   UND1 : ND2_654 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_653 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_652 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_217 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_217;

architecture SYN_STRUCTURAL of MUX21_217 is

   component ND2_649
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_650
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_651
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_217
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_217 port map( A => S, Y => SB);
   UND1 : ND2_651 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_650 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_649 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_216 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_216;

architecture SYN_STRUCTURAL of MUX21_216 is

   component ND2_646
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_647
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_648
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_216
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_216 port map( A => S, Y => SB);
   UND1 : ND2_648 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_647 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_646 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_215 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_215;

architecture SYN_STRUCTURAL of MUX21_215 is

   component ND2_643
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_644
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_645
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_215
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_215 port map( A => S, Y => SB);
   UND1 : ND2_645 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_644 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_643 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_214 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_214;

architecture SYN_STRUCTURAL of MUX21_214 is

   component ND2_640
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_641
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_642
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_214
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_214 port map( A => S, Y => SB);
   UND1 : ND2_642 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_641 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_640 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_213 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_213;

architecture SYN_STRUCTURAL of MUX21_213 is

   component ND2_637
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_638
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_639
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_213
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_213 port map( A => S, Y => SB);
   UND1 : ND2_639 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_638 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_637 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_212 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_212;

architecture SYN_STRUCTURAL of MUX21_212 is

   component ND2_634
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_635
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_636
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_212
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_212 port map( A => S, Y => SB);
   UND1 : ND2_636 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_635 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_634 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_211 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_211;

architecture SYN_STRUCTURAL of MUX21_211 is

   component ND2_631
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_632
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_633
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_211
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_211 port map( A => S, Y => SB);
   UND1 : ND2_633 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_632 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_631 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_210 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_210;

architecture SYN_STRUCTURAL of MUX21_210 is

   component ND2_628
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_629
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_630
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_210
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_210 port map( A => S, Y => SB);
   UND1 : ND2_630 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_629 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_628 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_209 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_209;

architecture SYN_STRUCTURAL of MUX21_209 is

   component ND2_625
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_626
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_627
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_209
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_209 port map( A => S, Y => SB);
   UND1 : ND2_627 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_626 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_625 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_208 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_208;

architecture SYN_STRUCTURAL of MUX21_208 is

   component ND2_622
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_623
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_624
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_208
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_208 port map( A => S, Y => SB);
   UND1 : ND2_624 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_623 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_622 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_207 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_207;

architecture SYN_STRUCTURAL of MUX21_207 is

   component ND2_619
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_620
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_621
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_207
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_207 port map( A => S, Y => SB);
   UND1 : ND2_621 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_620 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_619 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_206 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_206;

architecture SYN_STRUCTURAL of MUX21_206 is

   component ND2_616
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_617
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_618
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_206
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_206 port map( A => S, Y => SB);
   UND1 : ND2_618 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_617 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_616 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_205 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_205;

architecture SYN_STRUCTURAL of MUX21_205 is

   component ND2_613
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_614
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_615
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_205
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_205 port map( A => S, Y => SB);
   UND1 : ND2_615 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_614 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_613 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_204 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_204;

architecture SYN_STRUCTURAL of MUX21_204 is

   component ND2_610
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_611
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_612
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_204
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_204 port map( A => S, Y => SB);
   UND1 : ND2_612 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_611 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_610 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_203 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_203;

architecture SYN_STRUCTURAL of MUX21_203 is

   component ND2_607
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_608
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_609
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_203
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_203 port map( A => S, Y => SB);
   UND1 : ND2_609 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_608 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_607 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_202 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_202;

architecture SYN_STRUCTURAL of MUX21_202 is

   component ND2_604
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_605
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_606
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_202
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_202 port map( A => S, Y => SB);
   UND1 : ND2_606 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_605 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_604 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_201 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_201;

architecture SYN_STRUCTURAL of MUX21_201 is

   component ND2_601
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_602
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_603
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_201
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_201 port map( A => S, Y => SB);
   UND1 : ND2_603 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_602 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_601 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_200 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_200;

architecture SYN_STRUCTURAL of MUX21_200 is

   component ND2_598
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_599
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_600
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_200
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_200 port map( A => S, Y => SB);
   UND1 : ND2_600 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_599 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_598 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_199 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_199;

architecture SYN_STRUCTURAL of MUX21_199 is

   component ND2_595
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_596
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_597
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_199
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_199 port map( A => S, Y => SB);
   UND1 : ND2_597 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_596 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_595 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_198 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_198;

architecture SYN_STRUCTURAL of MUX21_198 is

   component ND2_592
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_593
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_594
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_198
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_198 port map( A => S, Y => SB);
   UND1 : ND2_594 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_593 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_592 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_197 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_197;

architecture SYN_STRUCTURAL of MUX21_197 is

   component ND2_589
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_590
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_591
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_197
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_197 port map( A => S, Y => SB);
   UND1 : ND2_591 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_590 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_589 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_196 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_196;

architecture SYN_STRUCTURAL of MUX21_196 is

   component ND2_586
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_587
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_588
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_196
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_196 port map( A => S, Y => SB);
   UND1 : ND2_588 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_587 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_586 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_195 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_195;

architecture SYN_STRUCTURAL of MUX21_195 is

   component ND2_583
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_584
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_585
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_195
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_195 port map( A => S, Y => SB);
   UND1 : ND2_585 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_584 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_583 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_194 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_194;

architecture SYN_STRUCTURAL of MUX21_194 is

   component ND2_580
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_581
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_582
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_194
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_194 port map( A => S, Y => SB);
   UND1 : ND2_582 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_581 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_580 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_193 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_193;

architecture SYN_STRUCTURAL of MUX21_193 is

   component ND2_577
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_578
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_579
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_193
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_193 port map( A => S, Y => SB);
   UND1 : ND2_579 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_578 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_577 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_192 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_192;

architecture SYN_STRUCTURAL of MUX21_192 is

   component ND2_574
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_575
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_576
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_192
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_192 port map( A => S, Y => SB);
   UND1 : ND2_576 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_575 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_574 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_191 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_191;

architecture SYN_STRUCTURAL of MUX21_191 is

   component ND2_571
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_572
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_573
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_191
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_191 port map( A => S, Y => SB);
   UND1 : ND2_573 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_572 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_571 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_190 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_190;

architecture SYN_STRUCTURAL of MUX21_190 is

   component ND2_568
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_569
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_570
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_190
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_190 port map( A => S, Y => SB);
   UND1 : ND2_570 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_569 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_568 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_189 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_189;

architecture SYN_STRUCTURAL of MUX21_189 is

   component ND2_565
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_566
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_567
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_189
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_189 port map( A => S, Y => SB);
   UND1 : ND2_567 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_566 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_565 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_188 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_188;

architecture SYN_STRUCTURAL of MUX21_188 is

   component ND2_562
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_563
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_564
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_188
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_188 port map( A => S, Y => SB);
   UND1 : ND2_564 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_563 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_562 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_187 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_187;

architecture SYN_STRUCTURAL of MUX21_187 is

   component ND2_559
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_560
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_561
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_187
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_187 port map( A => S, Y => SB);
   UND1 : ND2_561 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_560 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_559 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_186 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_186;

architecture SYN_STRUCTURAL of MUX21_186 is

   component ND2_556
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_557
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_558
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_186
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_186 port map( A => S, Y => SB);
   UND1 : ND2_558 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_557 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_556 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_185 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_185;

architecture SYN_STRUCTURAL of MUX21_185 is

   component ND2_553
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_554
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_555
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_185
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_185 port map( A => S, Y => SB);
   UND1 : ND2_555 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_554 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_553 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_184 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_184;

architecture SYN_STRUCTURAL of MUX21_184 is

   component ND2_550
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_551
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_552
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_184
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_184 port map( A => S, Y => SB);
   UND1 : ND2_552 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_551 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_550 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_183 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_183;

architecture SYN_STRUCTURAL of MUX21_183 is

   component ND2_547
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_548
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_549
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_183
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_183 port map( A => S, Y => SB);
   UND1 : ND2_549 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_548 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_547 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_182 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_182;

architecture SYN_STRUCTURAL of MUX21_182 is

   component ND2_544
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_545
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_546
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_182
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_182 port map( A => S, Y => SB);
   UND1 : ND2_546 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_545 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_544 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_181 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_181;

architecture SYN_STRUCTURAL of MUX21_181 is

   component ND2_541
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_542
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_543
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_181
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_181 port map( A => S, Y => SB);
   UND1 : ND2_543 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_542 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_541 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_180 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_180;

architecture SYN_STRUCTURAL of MUX21_180 is

   component ND2_538
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_539
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_540
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_180
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_180 port map( A => S, Y => SB);
   UND1 : ND2_540 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_539 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_538 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_179 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_179;

architecture SYN_STRUCTURAL of MUX21_179 is

   component ND2_535
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_536
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_537
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_179
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_179 port map( A => S, Y => SB);
   UND1 : ND2_537 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_536 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_535 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_178 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_178;

architecture SYN_STRUCTURAL of MUX21_178 is

   component ND2_532
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_533
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_534
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_178
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_178 port map( A => S, Y => SB);
   UND1 : ND2_534 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_533 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_532 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_177 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_177;

architecture SYN_STRUCTURAL of MUX21_177 is

   component ND2_529
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_530
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_531
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_177
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_177 port map( A => S, Y => SB);
   UND1 : ND2_531 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_530 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_529 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_176 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_176;

architecture SYN_STRUCTURAL of MUX21_176 is

   component ND2_526
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_527
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_528
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_176
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_176 port map( A => S, Y => SB);
   UND1 : ND2_528 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_527 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_526 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_175 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_175;

architecture SYN_STRUCTURAL of MUX21_175 is

   component ND2_523
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_524
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_525
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_175
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_175 port map( A => S, Y => SB);
   UND1 : ND2_525 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_524 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_523 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_174 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_174;

architecture SYN_STRUCTURAL of MUX21_174 is

   component ND2_520
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_521
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_522
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_174
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_174 port map( A => S, Y => SB);
   UND1 : ND2_522 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_521 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_520 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_173 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_173;

architecture SYN_STRUCTURAL of MUX21_173 is

   component ND2_517
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_518
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_519
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_173
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_173 port map( A => S, Y => SB);
   UND1 : ND2_519 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_518 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_517 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_172 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_172;

architecture SYN_STRUCTURAL of MUX21_172 is

   component ND2_514
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_515
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_516
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_172
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_172 port map( A => S, Y => SB);
   UND1 : ND2_516 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_515 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_514 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_171 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_171;

architecture SYN_STRUCTURAL of MUX21_171 is

   component ND2_511
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_512
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_513
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_171
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_171 port map( A => S, Y => SB);
   UND1 : ND2_513 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_512 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_511 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_170 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_170;

architecture SYN_STRUCTURAL of MUX21_170 is

   component ND2_508
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_509
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_510
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_170
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_170 port map( A => S, Y => SB);
   UND1 : ND2_510 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_509 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_508 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_169 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_169;

architecture SYN_STRUCTURAL of MUX21_169 is

   component ND2_505
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_506
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_507
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_169
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_169 port map( A => S, Y => SB);
   UND1 : ND2_507 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_506 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_505 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_168 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_168;

architecture SYN_STRUCTURAL of MUX21_168 is

   component ND2_502
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_503
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_504
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_168
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_168 port map( A => S, Y => SB);
   UND1 : ND2_504 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_503 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_502 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_167 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_167;

architecture SYN_STRUCTURAL of MUX21_167 is

   component ND2_499
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_500
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_501
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_167
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_167 port map( A => S, Y => SB);
   UND1 : ND2_501 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_500 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_499 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_166 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_166;

architecture SYN_STRUCTURAL of MUX21_166 is

   component ND2_496
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_497
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_498
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_166
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_166 port map( A => S, Y => SB);
   UND1 : ND2_498 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_497 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_496 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_165 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_165;

architecture SYN_STRUCTURAL of MUX21_165 is

   component ND2_493
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_494
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_495
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_165
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_165 port map( A => S, Y => SB);
   UND1 : ND2_495 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_494 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_493 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_164 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_164;

architecture SYN_STRUCTURAL of MUX21_164 is

   component ND2_490
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_491
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_492
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_164
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_164 port map( A => S, Y => SB);
   UND1 : ND2_492 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_491 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_490 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_163 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_163;

architecture SYN_STRUCTURAL of MUX21_163 is

   component ND2_487
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_488
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_489
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_163
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_163 port map( A => S, Y => SB);
   UND1 : ND2_489 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_488 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_487 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_162 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_162;

architecture SYN_STRUCTURAL of MUX21_162 is

   component ND2_484
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_485
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_486
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_162
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_162 port map( A => S, Y => SB);
   UND1 : ND2_486 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_485 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_484 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_161 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_161;

architecture SYN_STRUCTURAL of MUX21_161 is

   component ND2_481
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_482
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_483
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_161
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_161 port map( A => S, Y => SB);
   UND1 : ND2_483 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_482 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_481 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_160 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_160;

architecture SYN_STRUCTURAL of MUX21_160 is

   component ND2_478
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_479
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_480
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_160
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_160 port map( A => S, Y => SB);
   UND1 : ND2_480 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_479 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_478 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_159 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_159;

architecture SYN_STRUCTURAL of MUX21_159 is

   component ND2_475
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_476
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_477
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_159
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_159 port map( A => S, Y => SB);
   UND1 : ND2_477 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_476 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_475 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_158 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_158;

architecture SYN_STRUCTURAL of MUX21_158 is

   component ND2_472
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_473
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_474
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_158
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_158 port map( A => S, Y => SB);
   UND1 : ND2_474 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_473 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_472 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_157 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_157;

architecture SYN_STRUCTURAL of MUX21_157 is

   component ND2_469
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_470
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_471
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_157
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_157 port map( A => S, Y => SB);
   UND1 : ND2_471 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_470 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_469 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_156 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_156;

architecture SYN_STRUCTURAL of MUX21_156 is

   component ND2_466
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_467
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_468
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_156
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_156 port map( A => S, Y => SB);
   UND1 : ND2_468 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_467 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_466 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_155 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_155;

architecture SYN_STRUCTURAL of MUX21_155 is

   component ND2_463
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_464
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_465
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_155
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_155 port map( A => S, Y => SB);
   UND1 : ND2_465 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_464 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_463 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_154 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_154;

architecture SYN_STRUCTURAL of MUX21_154 is

   component ND2_460
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_461
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_462
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_154
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_154 port map( A => S, Y => SB);
   UND1 : ND2_462 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_461 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_460 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_153 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_153;

architecture SYN_STRUCTURAL of MUX21_153 is

   component ND2_457
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_458
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_459
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_153
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_153 port map( A => S, Y => SB);
   UND1 : ND2_459 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_458 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_457 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_152 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_152;

architecture SYN_STRUCTURAL of MUX21_152 is

   component ND2_454
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_455
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_456
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_152
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_152 port map( A => S, Y => SB);
   UND1 : ND2_456 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_455 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_454 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_151 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_151;

architecture SYN_STRUCTURAL of MUX21_151 is

   component ND2_451
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_452
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_453
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_151
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_151 port map( A => S, Y => SB);
   UND1 : ND2_453 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_452 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_451 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_150 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_150;

architecture SYN_STRUCTURAL of MUX21_150 is

   component ND2_448
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_449
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_450
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_150
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_150 port map( A => S, Y => SB);
   UND1 : ND2_450 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_449 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_448 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_149 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_149;

architecture SYN_STRUCTURAL of MUX21_149 is

   component ND2_445
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_446
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_447
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_149
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_149 port map( A => S, Y => SB);
   UND1 : ND2_447 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_446 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_445 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_148 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_148;

architecture SYN_STRUCTURAL of MUX21_148 is

   component ND2_442
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_443
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_444
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_148
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_148 port map( A => S, Y => SB);
   UND1 : ND2_444 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_443 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_442 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_147 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_147;

architecture SYN_STRUCTURAL of MUX21_147 is

   component ND2_439
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_440
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_441
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_147
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_147 port map( A => S, Y => SB);
   UND1 : ND2_441 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_440 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_439 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_146 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_146;

architecture SYN_STRUCTURAL of MUX21_146 is

   component ND2_436
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_437
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_438
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_146
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_146 port map( A => S, Y => SB);
   UND1 : ND2_438 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_437 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_436 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_145 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_145;

architecture SYN_STRUCTURAL of MUX21_145 is

   component ND2_433
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_434
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_435
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_145
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_145 port map( A => S, Y => SB);
   UND1 : ND2_435 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_434 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_433 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_144 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_144;

architecture SYN_STRUCTURAL of MUX21_144 is

   component ND2_430
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_431
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_432
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_144
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_144 port map( A => S, Y => SB);
   UND1 : ND2_432 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_431 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_430 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_143 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_143;

architecture SYN_STRUCTURAL of MUX21_143 is

   component ND2_427
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_428
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_429
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_143
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_143 port map( A => S, Y => SB);
   UND1 : ND2_429 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_428 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_427 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_142 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_142;

architecture SYN_STRUCTURAL of MUX21_142 is

   component ND2_424
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_425
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_426
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_142
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_142 port map( A => S, Y => SB);
   UND1 : ND2_426 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_425 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_424 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_141 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_141;

architecture SYN_STRUCTURAL of MUX21_141 is

   component ND2_421
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_422
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_423
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_141
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_141 port map( A => S, Y => SB);
   UND1 : ND2_423 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_422 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_421 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_140 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_140;

architecture SYN_STRUCTURAL of MUX21_140 is

   component ND2_418
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_419
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_420
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_140
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_140 port map( A => S, Y => SB);
   UND1 : ND2_420 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_419 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_418 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_139 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_139;

architecture SYN_STRUCTURAL of MUX21_139 is

   component ND2_415
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_416
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_417
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_139
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_139 port map( A => S, Y => SB);
   UND1 : ND2_417 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_416 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_415 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_138 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_138;

architecture SYN_STRUCTURAL of MUX21_138 is

   component ND2_412
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_413
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_414
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_138
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_138 port map( A => S, Y => SB);
   UND1 : ND2_414 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_413 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_412 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_137 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_137;

architecture SYN_STRUCTURAL of MUX21_137 is

   component ND2_409
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_410
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_411
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_137
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_137 port map( A => S, Y => SB);
   UND1 : ND2_411 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_410 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_409 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_136 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_136;

architecture SYN_STRUCTURAL of MUX21_136 is

   component ND2_406
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_407
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_408
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_136
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_136 port map( A => S, Y => SB);
   UND1 : ND2_408 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_407 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_406 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_135 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_135;

architecture SYN_STRUCTURAL of MUX21_135 is

   component ND2_403
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_404
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_405
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_135
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_135 port map( A => S, Y => SB);
   UND1 : ND2_405 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_404 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_403 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_134 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_134;

architecture SYN_STRUCTURAL of MUX21_134 is

   component ND2_400
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_401
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_402
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_134
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_134 port map( A => S, Y => SB);
   UND1 : ND2_402 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_401 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_400 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_133 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_133;

architecture SYN_STRUCTURAL of MUX21_133 is

   component ND2_397
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_398
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_399
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_133
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_133 port map( A => S, Y => SB);
   UND1 : ND2_399 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_398 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_397 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_132 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_132;

architecture SYN_STRUCTURAL of MUX21_132 is

   component ND2_394
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_395
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_396
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_132
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_132 port map( A => S, Y => SB);
   UND1 : ND2_396 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_395 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_394 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_131 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_131;

architecture SYN_STRUCTURAL of MUX21_131 is

   component ND2_391
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_392
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_393
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_131
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_131 port map( A => S, Y => SB);
   UND1 : ND2_393 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_392 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_391 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_130 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_130;

architecture SYN_STRUCTURAL of MUX21_130 is

   component ND2_388
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_389
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_390
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_130
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_130 port map( A => S, Y => SB);
   UND1 : ND2_390 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_389 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_388 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_129 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_129;

architecture SYN_STRUCTURAL of MUX21_129 is

   component ND2_385
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_386
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_387
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_129
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_129 port map( A => S, Y => SB);
   UND1 : ND2_387 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_386 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_385 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_128 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_128;

architecture SYN_STRUCTURAL of MUX21_128 is

   component ND2_382
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_383
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_384
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_128
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_128 port map( A => S, Y => SB);
   UND1 : ND2_384 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_383 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_382 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_127 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_127;

architecture SYN_STRUCTURAL of MUX21_127 is

   component ND2_379
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_380
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_381
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_127
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_127 port map( A => S, Y => SB);
   UND1 : ND2_381 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_380 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_379 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_126 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_126;

architecture SYN_STRUCTURAL of MUX21_126 is

   component ND2_376
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_377
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_378
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_126
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_126 port map( A => S, Y => SB);
   UND1 : ND2_378 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_377 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_376 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_125 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_125;

architecture SYN_STRUCTURAL of MUX21_125 is

   component ND2_373
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_374
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_375
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_125
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_125 port map( A => S, Y => SB);
   UND1 : ND2_375 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_374 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_373 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_124 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_124;

architecture SYN_STRUCTURAL of MUX21_124 is

   component ND2_370
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_371
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_372
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_124
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_124 port map( A => S, Y => SB);
   UND1 : ND2_372 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_371 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_370 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_123 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_123;

architecture SYN_STRUCTURAL of MUX21_123 is

   component ND2_367
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_368
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_369
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_123
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_123 port map( A => S, Y => SB);
   UND1 : ND2_369 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_368 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_367 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_122 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_122;

architecture SYN_STRUCTURAL of MUX21_122 is

   component ND2_364
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_365
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_366
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_122
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_122 port map( A => S, Y => SB);
   UND1 : ND2_366 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_365 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_364 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_121 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_121;

architecture SYN_STRUCTURAL of MUX21_121 is

   component ND2_361
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_362
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_363
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_121
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_121 port map( A => S, Y => SB);
   UND1 : ND2_363 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_362 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_361 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_120 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_120;

architecture SYN_STRUCTURAL of MUX21_120 is

   component ND2_358
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_359
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_360
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_120
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_120 port map( A => S, Y => SB);
   UND1 : ND2_360 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_359 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_358 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_119 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_119;

architecture SYN_STRUCTURAL of MUX21_119 is

   component ND2_355
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_356
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_357
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_119
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_119 port map( A => S, Y => SB);
   UND1 : ND2_357 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_356 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_355 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_118 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_118;

architecture SYN_STRUCTURAL of MUX21_118 is

   component ND2_352
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_353
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_354
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_118
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_118 port map( A => S, Y => SB);
   UND1 : ND2_354 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_353 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_352 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_117 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_117;

architecture SYN_STRUCTURAL of MUX21_117 is

   component ND2_349
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_350
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_351
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_117
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_117 port map( A => S, Y => SB);
   UND1 : ND2_351 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_350 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_349 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_116 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_116;

architecture SYN_STRUCTURAL of MUX21_116 is

   component ND2_346
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_347
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_348
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_116
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_116 port map( A => S, Y => SB);
   UND1 : ND2_348 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_347 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_346 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_115 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_115;

architecture SYN_STRUCTURAL of MUX21_115 is

   component ND2_343
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_344
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_345
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_115
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_115 port map( A => S, Y => SB);
   UND1 : ND2_345 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_344 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_343 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_114 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_114;

architecture SYN_STRUCTURAL of MUX21_114 is

   component ND2_340
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_341
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_342
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_114
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_114 port map( A => S, Y => SB);
   UND1 : ND2_342 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_341 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_340 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_113 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_113;

architecture SYN_STRUCTURAL of MUX21_113 is

   component ND2_337
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_338
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_339
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_113
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_113 port map( A => S, Y => SB);
   UND1 : ND2_339 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_338 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_337 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_112 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_112;

architecture SYN_STRUCTURAL of MUX21_112 is

   component ND2_334
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_335
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_336
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_112
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_112 port map( A => S, Y => SB);
   UND1 : ND2_336 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_335 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_334 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_111 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_111;

architecture SYN_STRUCTURAL of MUX21_111 is

   component ND2_331
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_332
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_333
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_111
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_111 port map( A => S, Y => SB);
   UND1 : ND2_333 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_332 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_331 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_110 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_110;

architecture SYN_STRUCTURAL of MUX21_110 is

   component ND2_328
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_329
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_330
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_110
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_110 port map( A => S, Y => SB);
   UND1 : ND2_330 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_329 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_328 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_109 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_109;

architecture SYN_STRUCTURAL of MUX21_109 is

   component ND2_325
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_326
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_327
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_109
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_109 port map( A => S, Y => SB);
   UND1 : ND2_327 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_326 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_325 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_108 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_108;

architecture SYN_STRUCTURAL of MUX21_108 is

   component ND2_322
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_323
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_324
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_108
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_108 port map( A => S, Y => SB);
   UND1 : ND2_324 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_323 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_322 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_107 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_107;

architecture SYN_STRUCTURAL of MUX21_107 is

   component ND2_319
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_320
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_321
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_107
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_107 port map( A => S, Y => SB);
   UND1 : ND2_321 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_320 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_319 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_106 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_106;

architecture SYN_STRUCTURAL of MUX21_106 is

   component ND2_316
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_317
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_318
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_106
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_106 port map( A => S, Y => SB);
   UND1 : ND2_318 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_317 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_316 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_105 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_105;

architecture SYN_STRUCTURAL of MUX21_105 is

   component ND2_313
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_314
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_315
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_105
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_105 port map( A => S, Y => SB);
   UND1 : ND2_315 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_314 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_313 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_104 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_104;

architecture SYN_STRUCTURAL of MUX21_104 is

   component ND2_310
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_311
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_312
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_104
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_104 port map( A => S, Y => SB);
   UND1 : ND2_312 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_311 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_310 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_103 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_103;

architecture SYN_STRUCTURAL of MUX21_103 is

   component ND2_307
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_308
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_309
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_103
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_103 port map( A => S, Y => SB);
   UND1 : ND2_309 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_308 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_307 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_102 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_102;

architecture SYN_STRUCTURAL of MUX21_102 is

   component ND2_304
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_305
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_306
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_102
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_102 port map( A => S, Y => SB);
   UND1 : ND2_306 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_305 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_304 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_101 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_101;

architecture SYN_STRUCTURAL of MUX21_101 is

   component ND2_301
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_302
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_303
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_101
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_101 port map( A => S, Y => SB);
   UND1 : ND2_303 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_302 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_301 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_100 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_100;

architecture SYN_STRUCTURAL of MUX21_100 is

   component ND2_298
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_299
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_300
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_100
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_100 port map( A => S, Y => SB);
   UND1 : ND2_300 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_299 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_298 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_99 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_99;

architecture SYN_STRUCTURAL of MUX21_99 is

   component ND2_295
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_296
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_297
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_99
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_99 port map( A => S, Y => SB);
   UND1 : ND2_297 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_296 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_295 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_98 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_98;

architecture SYN_STRUCTURAL of MUX21_98 is

   component ND2_292
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_293
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_294
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_98
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_98 port map( A => S, Y => SB);
   UND1 : ND2_294 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_293 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_292 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_97 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_97;

architecture SYN_STRUCTURAL of MUX21_97 is

   component ND2_289
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_290
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_291
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_97
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_97 port map( A => S, Y => SB);
   UND1 : ND2_291 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_290 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_289 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_96 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_96;

architecture SYN_STRUCTURAL of MUX21_96 is

   component ND2_286
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_287
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_288
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_96
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_96 port map( A => S, Y => SB);
   UND1 : ND2_288 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_287 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_286 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_95 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_95;

architecture SYN_STRUCTURAL of MUX21_95 is

   component ND2_283
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_284
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_285
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_95
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_95 port map( A => S, Y => SB);
   UND1 : ND2_285 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_284 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_283 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_94 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_94;

architecture SYN_STRUCTURAL of MUX21_94 is

   component ND2_280
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_281
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_282
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_94
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_94 port map( A => S, Y => SB);
   UND1 : ND2_282 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_281 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_280 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_93 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_93;

architecture SYN_STRUCTURAL of MUX21_93 is

   component ND2_277
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_278
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_279
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_93
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_93 port map( A => S, Y => SB);
   UND1 : ND2_279 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_278 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_277 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_92 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_92;

architecture SYN_STRUCTURAL of MUX21_92 is

   component ND2_274
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_275
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_276
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_92
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_92 port map( A => S, Y => SB);
   UND1 : ND2_276 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_275 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_274 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_91 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_91;

architecture SYN_STRUCTURAL of MUX21_91 is

   component ND2_271
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_272
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_273
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_91
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_91 port map( A => S, Y => SB);
   UND1 : ND2_273 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_272 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_271 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_90 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_90;

architecture SYN_STRUCTURAL of MUX21_90 is

   component ND2_268
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_269
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_270
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_90
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_90 port map( A => S, Y => SB);
   UND1 : ND2_270 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_269 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_268 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_89 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_89;

architecture SYN_STRUCTURAL of MUX21_89 is

   component ND2_265
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_266
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_267
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_89
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_89 port map( A => S, Y => SB);
   UND1 : ND2_267 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_266 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_265 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_88 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_88;

architecture SYN_STRUCTURAL of MUX21_88 is

   component ND2_262
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_263
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_264
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_88
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_88 port map( A => S, Y => SB);
   UND1 : ND2_264 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_263 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_262 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_87 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_87;

architecture SYN_STRUCTURAL of MUX21_87 is

   component ND2_259
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_260
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_261
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_87
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_87 port map( A => S, Y => SB);
   UND1 : ND2_261 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_260 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_259 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_86 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_86;

architecture SYN_STRUCTURAL of MUX21_86 is

   component ND2_256
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_257
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_258
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_86
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_86 port map( A => S, Y => SB);
   UND1 : ND2_258 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_257 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_256 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_85 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_85;

architecture SYN_STRUCTURAL of MUX21_85 is

   component ND2_253
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_254
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_255
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_85
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_85 port map( A => S, Y => SB);
   UND1 : ND2_255 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_254 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_253 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_84 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_84;

architecture SYN_STRUCTURAL of MUX21_84 is

   component ND2_250
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_251
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_252
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_84
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_84 port map( A => S, Y => SB);
   UND1 : ND2_252 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_251 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_250 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_83 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_83;

architecture SYN_STRUCTURAL of MUX21_83 is

   component ND2_247
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_248
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_249
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_83
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_83 port map( A => S, Y => SB);
   UND1 : ND2_249 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_248 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_247 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_82 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_82;

architecture SYN_STRUCTURAL of MUX21_82 is

   component ND2_244
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_245
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_246
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_82
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_82 port map( A => S, Y => SB);
   UND1 : ND2_246 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_245 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_244 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_81 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_81;

architecture SYN_STRUCTURAL of MUX21_81 is

   component ND2_241
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_242
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_243
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_81
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_81 port map( A => S, Y => SB);
   UND1 : ND2_243 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_242 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_241 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_80 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_80;

architecture SYN_STRUCTURAL of MUX21_80 is

   component ND2_238
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_239
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_240
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_80
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_80 port map( A => S, Y => SB);
   UND1 : ND2_240 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_239 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_238 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_79 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_79;

architecture SYN_STRUCTURAL of MUX21_79 is

   component ND2_235
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_236
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_237
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_79
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_79 port map( A => S, Y => SB);
   UND1 : ND2_237 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_236 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_235 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_78 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_78;

architecture SYN_STRUCTURAL of MUX21_78 is

   component ND2_232
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_233
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_234
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_78
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_78 port map( A => S, Y => SB);
   UND1 : ND2_234 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_233 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_232 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_77 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_77;

architecture SYN_STRUCTURAL of MUX21_77 is

   component ND2_229
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_230
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_231
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_77
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_77 port map( A => S, Y => SB);
   UND1 : ND2_231 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_230 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_229 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_76 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_76;

architecture SYN_STRUCTURAL of MUX21_76 is

   component ND2_226
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_227
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_228
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_76
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_76 port map( A => S, Y => SB);
   UND1 : ND2_228 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_227 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_226 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_75 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_75;

architecture SYN_STRUCTURAL of MUX21_75 is

   component ND2_223
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_224
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_225
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_75
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_75 port map( A => S, Y => SB);
   UND1 : ND2_225 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_224 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_223 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_74 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_74;

architecture SYN_STRUCTURAL of MUX21_74 is

   component ND2_220
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_221
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_222
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_74
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_74 port map( A => S, Y => SB);
   UND1 : ND2_222 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_221 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_220 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_73 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_73;

architecture SYN_STRUCTURAL of MUX21_73 is

   component ND2_217
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_218
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_219
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_73
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_73 port map( A => S, Y => SB);
   UND1 : ND2_219 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_218 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_217 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_72 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_72;

architecture SYN_STRUCTURAL of MUX21_72 is

   component ND2_214
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_215
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_216
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_72
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_72 port map( A => S, Y => SB);
   UND1 : ND2_216 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_215 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_214 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_71 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_71;

architecture SYN_STRUCTURAL of MUX21_71 is

   component ND2_211
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_212
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_213
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_71
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_71 port map( A => S, Y => SB);
   UND1 : ND2_213 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_212 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_211 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_70 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_70;

architecture SYN_STRUCTURAL of MUX21_70 is

   component ND2_208
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_209
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_210
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_70
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_70 port map( A => S, Y => SB);
   UND1 : ND2_210 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_209 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_208 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_69 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_69;

architecture SYN_STRUCTURAL of MUX21_69 is

   component ND2_205
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_206
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_207
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_69
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_69 port map( A => S, Y => SB);
   UND1 : ND2_207 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_206 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_205 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_68 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_68;

architecture SYN_STRUCTURAL of MUX21_68 is

   component ND2_202
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_203
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_204
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_68
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_68 port map( A => S, Y => SB);
   UND1 : ND2_204 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_203 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_202 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_67 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_67;

architecture SYN_STRUCTURAL of MUX21_67 is

   component ND2_199
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_200
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_201
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_67
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_67 port map( A => S, Y => SB);
   UND1 : ND2_201 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_200 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_199 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_66 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_66;

architecture SYN_STRUCTURAL of MUX21_66 is

   component ND2_196
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_197
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_198
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_66
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_66 port map( A => S, Y => SB);
   UND1 : ND2_198 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_197 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_196 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_65 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_65;

architecture SYN_STRUCTURAL of MUX21_65 is

   component ND2_193
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_194
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_195
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_65
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_65 port map( A => S, Y => SB);
   UND1 : ND2_195 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_194 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_193 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_64 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_64;

architecture SYN_STRUCTURAL of MUX21_64 is

   component ND2_190
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_191
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_192
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_64
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_64 port map( A => S, Y => SB);
   UND1 : ND2_192 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_191 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_190 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_63 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_63;

architecture SYN_STRUCTURAL of MUX21_63 is

   component ND2_187
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_188
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_189
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_63
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_63 port map( A => S, Y => SB);
   UND1 : ND2_189 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_188 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_187 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_62 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_62;

architecture SYN_STRUCTURAL of MUX21_62 is

   component ND2_184
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_185
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_186
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_62
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_62 port map( A => S, Y => SB);
   UND1 : ND2_186 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_185 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_184 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_61 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_61;

architecture SYN_STRUCTURAL of MUX21_61 is

   component ND2_181
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_182
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_183
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_61
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_61 port map( A => S, Y => SB);
   UND1 : ND2_183 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_182 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_181 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_60 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_60;

architecture SYN_STRUCTURAL of MUX21_60 is

   component ND2_178
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_179
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_180
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_60
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_60 port map( A => S, Y => SB);
   UND1 : ND2_180 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_179 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_178 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_59 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_59;

architecture SYN_STRUCTURAL of MUX21_59 is

   component ND2_175
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_176
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_177
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_59
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_59 port map( A => S, Y => SB);
   UND1 : ND2_177 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_176 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_175 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_58 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_58;

architecture SYN_STRUCTURAL of MUX21_58 is

   component ND2_172
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_173
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_174
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_58
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_58 port map( A => S, Y => SB);
   UND1 : ND2_174 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_173 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_172 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_57 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_57;

architecture SYN_STRUCTURAL of MUX21_57 is

   component ND2_169
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_170
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_171
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_57
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_57 port map( A => S, Y => SB);
   UND1 : ND2_171 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_170 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_169 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_56 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_56;

architecture SYN_STRUCTURAL of MUX21_56 is

   component ND2_166
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_167
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_168
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_56
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_56 port map( A => S, Y => SB);
   UND1 : ND2_168 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_167 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_166 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_55 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_55;

architecture SYN_STRUCTURAL of MUX21_55 is

   component ND2_163
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_164
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_165
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_55
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_55 port map( A => S, Y => SB);
   UND1 : ND2_165 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_164 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_163 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_54 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_54;

architecture SYN_STRUCTURAL of MUX21_54 is

   component ND2_160
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_161
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_162
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_54
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_54 port map( A => S, Y => SB);
   UND1 : ND2_162 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_161 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_160 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_53 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_53;

architecture SYN_STRUCTURAL of MUX21_53 is

   component ND2_157
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_158
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_159
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_53
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_53 port map( A => S, Y => SB);
   UND1 : ND2_159 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_158 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_157 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_52 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_52;

architecture SYN_STRUCTURAL of MUX21_52 is

   component ND2_154
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_155
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_156
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_52
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_52 port map( A => S, Y => SB);
   UND1 : ND2_156 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_155 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_154 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_51 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_51;

architecture SYN_STRUCTURAL of MUX21_51 is

   component ND2_151
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_152
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_153
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_51
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_51 port map( A => S, Y => SB);
   UND1 : ND2_153 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_152 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_151 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_50 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_50;

architecture SYN_STRUCTURAL of MUX21_50 is

   component ND2_148
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_149
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_150
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_50
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_50 port map( A => S, Y => SB);
   UND1 : ND2_150 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_149 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_148 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_49 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_49;

architecture SYN_STRUCTURAL of MUX21_49 is

   component ND2_145
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_146
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_147
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_49
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_49 port map( A => S, Y => SB);
   UND1 : ND2_147 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_146 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_145 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_48 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_48;

architecture SYN_STRUCTURAL of MUX21_48 is

   component ND2_142
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_143
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_144
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_48
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_48 port map( A => S, Y => SB);
   UND1 : ND2_144 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_143 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_142 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_47 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_47;

architecture SYN_STRUCTURAL of MUX21_47 is

   component ND2_139
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_140
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_141
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_47
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_47 port map( A => S, Y => SB);
   UND1 : ND2_141 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_140 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_139 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_46 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_46;

architecture SYN_STRUCTURAL of MUX21_46 is

   component ND2_136
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_137
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_138
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_46
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_46 port map( A => S, Y => SB);
   UND1 : ND2_138 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_137 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_136 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_45 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_45;

architecture SYN_STRUCTURAL of MUX21_45 is

   component ND2_133
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_134
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_135
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_45
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_45 port map( A => S, Y => SB);
   UND1 : ND2_135 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_134 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_133 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_44 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_44;

architecture SYN_STRUCTURAL of MUX21_44 is

   component ND2_130
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_131
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_132
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_44
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_44 port map( A => S, Y => SB);
   UND1 : ND2_132 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_131 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_130 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_43 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_43;

architecture SYN_STRUCTURAL of MUX21_43 is

   component ND2_127
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_128
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_129
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_43
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_43 port map( A => S, Y => SB);
   UND1 : ND2_129 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_128 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_127 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_42 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_42;

architecture SYN_STRUCTURAL of MUX21_42 is

   component ND2_124
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_125
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_126
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_42
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_42 port map( A => S, Y => SB);
   UND1 : ND2_126 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_125 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_124 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_41 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_41;

architecture SYN_STRUCTURAL of MUX21_41 is

   component ND2_121
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_122
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_123
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_41
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_41 port map( A => S, Y => SB);
   UND1 : ND2_123 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_122 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_121 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_40 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_40;

architecture SYN_STRUCTURAL of MUX21_40 is

   component ND2_118
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_119
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_120
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_40
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_40 port map( A => S, Y => SB);
   UND1 : ND2_120 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_119 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_118 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_39 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_39;

architecture SYN_STRUCTURAL of MUX21_39 is

   component ND2_115
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_116
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_117
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_39
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_39 port map( A => S, Y => SB);
   UND1 : ND2_117 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_116 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_115 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_38 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_38;

architecture SYN_STRUCTURAL of MUX21_38 is

   component ND2_112
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_113
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_114
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_38
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_38 port map( A => S, Y => SB);
   UND1 : ND2_114 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_113 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_112 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_37 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_37;

architecture SYN_STRUCTURAL of MUX21_37 is

   component ND2_109
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_110
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_111
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_37
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_37 port map( A => S, Y => SB);
   UND1 : ND2_111 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_110 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_109 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_36 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_36;

architecture SYN_STRUCTURAL of MUX21_36 is

   component ND2_106
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_107
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_108
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_36
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_36 port map( A => S, Y => SB);
   UND1 : ND2_108 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_107 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_106 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_35 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_35;

architecture SYN_STRUCTURAL of MUX21_35 is

   component ND2_103
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_104
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_105
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_35
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_35 port map( A => S, Y => SB);
   UND1 : ND2_105 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_104 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_103 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_34 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_34;

architecture SYN_STRUCTURAL of MUX21_34 is

   component ND2_100
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_101
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_102
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_34
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_34 port map( A => S, Y => SB);
   UND1 : ND2_102 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_101 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_100 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_33 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_33;

architecture SYN_STRUCTURAL of MUX21_33 is

   component ND2_97
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_98
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_99
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_33
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_33 port map( A => S, Y => SB);
   UND1 : ND2_99 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_98 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_97 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_32 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_32;

architecture SYN_STRUCTURAL of MUX21_32 is

   component ND2_94
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_95
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_96
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_32
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_32 port map( A => S, Y => SB);
   UND1 : ND2_96 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_95 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_94 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_31 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_31;

architecture SYN_STRUCTURAL of MUX21_31 is

   component ND2_91
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_92
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_93
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_31
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_31 port map( A => S, Y => SB);
   UND1 : ND2_93 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_92 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_91 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_30 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_30;

architecture SYN_STRUCTURAL of MUX21_30 is

   component ND2_88
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_89
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_90
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_30
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_30 port map( A => S, Y => SB);
   UND1 : ND2_90 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_89 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_88 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_29 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_29;

architecture SYN_STRUCTURAL of MUX21_29 is

   component ND2_85
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_86
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_87
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_29
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_29 port map( A => S, Y => SB);
   UND1 : ND2_87 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_86 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_85 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_28 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_28;

architecture SYN_STRUCTURAL of MUX21_28 is

   component ND2_82
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_83
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_84
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_28
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_28 port map( A => S, Y => SB);
   UND1 : ND2_84 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_83 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_82 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_27 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_27;

architecture SYN_STRUCTURAL_architecture of MUX21_27 is

   component ND2_79
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_80
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_81
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_27
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_27 port map( A => S, Y => SB);
   UND1 : ND2_81 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_80 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_79 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL_architecture;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_26 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_26;

architecture SYN_STRUCTURAL_architecture2 of MUX21_26 is

   component ND2_76
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_77
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_78
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_26
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_26 port map( A => S, Y => SB);
   UND1 : ND2_78 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_77 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_76 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL_architecture2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_25 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_25;

architecture SYN_STRUCTURAL_architecture3 of MUX21_25 is

   component ND2_73
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_74
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_75
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_25
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_25 port map( A => S, Y => SB);
   UND1 : ND2_75 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_74 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_73 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL_architecture3;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_24 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_24;

architecture SYN_STRUCTURAL of MUX21_24 is

   component ND2_70
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_71
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_72
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_24
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_24 port map( A => S, Y => SB);
   UND1 : ND2_72 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_71 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_70 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_23 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_23;

architecture SYN_STRUCTURAL_architecture of MUX21_23 is

   component ND2_67
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_68
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_69
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_23
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_23 port map( A => S, Y => SB);
   UND1 : ND2_69 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_68 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_67 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL_architecture;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_22 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_22;

architecture SYN_STRUCTURAL_architecture2 of MUX21_22 is

   component ND2_64
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_65
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_66
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_22
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_22 port map( A => S, Y => SB);
   UND1 : ND2_66 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_65 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_64 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL_architecture2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_21 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_21;

architecture SYN_STRUCTURAL_architecture3 of MUX21_21 is

   component ND2_61
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_62
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_63
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_21
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_21 port map( A => S, Y => SB);
   UND1 : ND2_63 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_62 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_61 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL_architecture3;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_20 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_20;

architecture SYN_STRUCTURAL of MUX21_20 is

   component ND2_58
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_59
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_60
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_20
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_20 port map( A => S, Y => SB);
   UND1 : ND2_60 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_59 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_58 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_19 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_19;

architecture SYN_STRUCTURAL_architecture of MUX21_19 is

   component ND2_55
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_56
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_57
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_19
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_19 port map( A => S, Y => SB);
   UND1 : ND2_57 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_56 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_55 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL_architecture;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_18 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_18;

architecture SYN_STRUCTURAL_architecture2 of MUX21_18 is

   component ND2_52
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_53
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_54
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_18
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_18 port map( A => S, Y => SB);
   UND1 : ND2_54 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_53 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_52 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL_architecture2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_17 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_17;

architecture SYN_STRUCTURAL_architecture3 of MUX21_17 is

   component ND2_49
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_50
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_51
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_17
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_17 port map( A => S, Y => SB);
   UND1 : ND2_51 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_50 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_49 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL_architecture3;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_16 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_16;

architecture SYN_STRUCTURAL of MUX21_16 is

   component ND2_46
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_47
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_48
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_16
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_16 port map( A => S, Y => SB);
   UND1 : ND2_48 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_47 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_46 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_15 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_15;

architecture SYN_STRUCTURAL_architecture of MUX21_15 is

   component ND2_43
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_44
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_45
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_15
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_15 port map( A => S, Y => SB);
   UND1 : ND2_45 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_44 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_43 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL_architecture;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_14 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_14;

architecture SYN_STRUCTURAL_architecture2 of MUX21_14 is

   component ND2_40
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_41
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_42
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_14
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_14 port map( A => S, Y => SB);
   UND1 : ND2_42 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_41 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_40 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL_architecture2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_13 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_13;

architecture SYN_STRUCTURAL_architecture3 of MUX21_13 is

   component ND2_37
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_38
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_39
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_13
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_13 port map( A => S, Y => SB);
   UND1 : ND2_39 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_38 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_37 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL_architecture3;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_12 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_12;

architecture SYN_STRUCTURAL of MUX21_12 is

   component ND2_34
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_35
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_36
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_12
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_12 port map( A => S, Y => SB);
   UND1 : ND2_36 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_35 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_34 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_11 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_11;

architecture SYN_STRUCTURAL_architecture of MUX21_11 is

   component ND2_31
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_32
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_33
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_11
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_11 port map( A => S, Y => SB);
   UND1 : ND2_33 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_32 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_31 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL_architecture;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_10 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_10;

architecture SYN_STRUCTURAL_architecture2 of MUX21_10 is

   component ND2_28
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_29
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_30
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_10
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_10 port map( A => S, Y => SB);
   UND1 : ND2_30 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_29 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_28 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL_architecture2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_9 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_9;

architecture SYN_STRUCTURAL_architecture3 of MUX21_9 is

   component ND2_25
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_26
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_27
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_9
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_9 port map( A => S, Y => SB);
   UND1 : ND2_27 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_26 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_25 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL_architecture3;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_8 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_8;

architecture SYN_STRUCTURAL of MUX21_8 is

   component ND2_22
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_23
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_24
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_8
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_8 port map( A => S, Y => SB);
   UND1 : ND2_24 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_23 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_22 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_7 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_7;

architecture SYN_STRUCTURAL_architecture of MUX21_7 is

   component ND2_19
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_20
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_21
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_7
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_7 port map( A => S, Y => SB);
   UND1 : ND2_21 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_20 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_19 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL_architecture;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_6 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_6;

architecture SYN_STRUCTURAL_architecture2 of MUX21_6 is

   component ND2_16
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_17
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_18
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_6
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_6 port map( A => S, Y => SB);
   UND1 : ND2_18 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_17 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_16 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL_architecture2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_5 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_5;

architecture SYN_STRUCTURAL_architecture3 of MUX21_5 is

   component ND2_13
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_14
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_15
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_5
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_5 port map( A => S, Y => SB);
   UND1 : ND2_15 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_14 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_13 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL_architecture3;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_4 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_4;

architecture SYN_STRUCTURAL of MUX21_4 is

   component ND2_10
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_11
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_12
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_4
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_4 port map( A => S, Y => SB);
   UND1 : ND2_12 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_11 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_10 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_3 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_3;

architecture SYN_STRUCTURAL_architecture of MUX21_3 is

   component ND2_7
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_8
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_9
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_3
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_3 port map( A => S, Y => SB);
   UND1 : ND2_9 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_8 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_7 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL_architecture;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_2 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_2;

architecture SYN_STRUCTURAL_architecture2 of MUX21_2 is

   component ND2_4
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_5
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_6
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_2
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_2 port map( A => S, Y => SB);
   UND1 : ND2_6 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_5 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_4 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL_architecture2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_1 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_1;

architecture SYN_STRUCTURAL_architecture3 of MUX21_1 is

   component ND2_1
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_2
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_3
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_1
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_1 port map( A => S, Y => SB);
   UND1 : ND2_3 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_2 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_1 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL_architecture3;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity regFFD_NBIT6_1 is

   port( CK, RESET, ENABLE : in std_logic;  D : in std_logic_vector (5 downto 
         0);  Q : out std_logic_vector (5 downto 0));

end regFFD_NBIT6_1;

architecture SYN_ASYNCHBEHAV of regFFD_NBIT6_1 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32,
      n33, n34, n35, n36 : std_logic;

begin
   
   Q_reg_5_inst : DFFR_X1 port map( D => n19, CK => CK, RN => RESET, Q => Q(5),
                           QN => n25);
   Q_reg_4_inst : DFFR_X1 port map( D => n20, CK => CK, RN => RESET, Q => Q(4),
                           QN => n26);
   Q_reg_3_inst : DFFR_X1 port map( D => n21, CK => CK, RN => RESET, Q => Q(3),
                           QN => n27);
   Q_reg_2_inst : DFFR_X1 port map( D => n22, CK => CK, RN => RESET, Q => Q(2),
                           QN => n28);
   Q_reg_1_inst : DFFR_X1 port map( D => n23, CK => CK, RN => RESET, Q => Q(1),
                           QN => n29);
   Q_reg_0_inst : DFFR_X1 port map( D => n24, CK => CK, RN => RESET, Q => Q(0),
                           QN => n30);
   U2 : OAI21_X1 port map( B1 => n30, B2 => ENABLE, A => n36, ZN => n24);
   U3 : NAND2_X1 port map( A1 => ENABLE, A2 => D(0), ZN => n36);
   U4 : OAI21_X1 port map( B1 => n29, B2 => ENABLE, A => n35, ZN => n23);
   U5 : NAND2_X1 port map( A1 => D(1), A2 => ENABLE, ZN => n35);
   U6 : OAI21_X1 port map( B1 => n28, B2 => ENABLE, A => n34, ZN => n22);
   U7 : NAND2_X1 port map( A1 => D(2), A2 => ENABLE, ZN => n34);
   U8 : OAI21_X1 port map( B1 => n27, B2 => ENABLE, A => n33, ZN => n21);
   U9 : NAND2_X1 port map( A1 => D(3), A2 => ENABLE, ZN => n33);
   U10 : OAI21_X1 port map( B1 => n26, B2 => ENABLE, A => n32, ZN => n20);
   U11 : NAND2_X1 port map( A1 => D(4), A2 => ENABLE, ZN => n32);
   U12 : OAI21_X1 port map( B1 => n25, B2 => ENABLE, A => n31, ZN => n19);
   U13 : NAND2_X1 port map( A1 => D(5), A2 => ENABLE, ZN => n31);

end SYN_ASYNCHBEHAV;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity regFFD_NBIT5_2 is

   port( CK, RESET, ENABLE : in std_logic;  D : in std_logic_vector (4 downto 
         0);  Q : out std_logic_vector (4 downto 0));

end regFFD_NBIT5_2;

architecture SYN_ASYNCHBEHAV of regFFD_NBIT5_2 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29,
      n30 : std_logic;

begin
   
   Q_reg_4_inst : DFFR_X1 port map( D => n16, CK => CK, RN => RESET, Q => Q(4),
                           QN => n21);
   Q_reg_3_inst : DFFR_X1 port map( D => n17, CK => CK, RN => RESET, Q => Q(3),
                           QN => n22);
   Q_reg_2_inst : DFFR_X1 port map( D => n18, CK => CK, RN => RESET, Q => Q(2),
                           QN => n23);
   Q_reg_1_inst : DFFR_X1 port map( D => n19, CK => CK, RN => RESET, Q => Q(1),
                           QN => n24);
   Q_reg_0_inst : DFFR_X1 port map( D => n20, CK => CK, RN => RESET, Q => Q(0),
                           QN => n25);
   U2 : OAI21_X1 port map( B1 => n25, B2 => ENABLE, A => n30, ZN => n20);
   U3 : NAND2_X1 port map( A1 => ENABLE, A2 => D(0), ZN => n30);
   U4 : OAI21_X1 port map( B1 => n24, B2 => ENABLE, A => n29, ZN => n19);
   U5 : NAND2_X1 port map( A1 => D(1), A2 => ENABLE, ZN => n29);
   U6 : OAI21_X1 port map( B1 => n23, B2 => ENABLE, A => n28, ZN => n18);
   U7 : NAND2_X1 port map( A1 => D(2), A2 => ENABLE, ZN => n28);
   U8 : OAI21_X1 port map( B1 => n22, B2 => ENABLE, A => n27, ZN => n17);
   U9 : NAND2_X1 port map( A1 => D(3), A2 => ENABLE, ZN => n27);
   U10 : OAI21_X1 port map( B1 => n21, B2 => ENABLE, A => n26, ZN => n16);
   U11 : NAND2_X1 port map( A1 => D(4), A2 => ENABLE, ZN => n26);

end SYN_ASYNCHBEHAV;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity regFFD_NBIT5_1 is

   port( CK, RESET, ENABLE : in std_logic;  D : in std_logic_vector (4 downto 
         0);  Q : out std_logic_vector (4 downto 0));

end regFFD_NBIT5_1;

architecture SYN_ASYNCHBEHAV of regFFD_NBIT5_1 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29,
      n30 : std_logic;

begin
   
   Q_reg_4_inst : DFFR_X1 port map( D => n16, CK => CK, RN => RESET, Q => Q(4),
                           QN => n21);
   Q_reg_3_inst : DFFR_X1 port map( D => n17, CK => CK, RN => RESET, Q => Q(3),
                           QN => n22);
   Q_reg_2_inst : DFFR_X1 port map( D => n18, CK => CK, RN => RESET, Q => Q(2),
                           QN => n23);
   Q_reg_1_inst : DFFR_X1 port map( D => n19, CK => CK, RN => RESET, Q => Q(1),
                           QN => n24);
   Q_reg_0_inst : DFFR_X1 port map( D => n20, CK => CK, RN => RESET, Q => Q(0),
                           QN => n25);
   U2 : OAI21_X1 port map( B1 => n25, B2 => ENABLE, A => n30, ZN => n20);
   U3 : NAND2_X1 port map( A1 => ENABLE, A2 => D(0), ZN => n30);
   U4 : OAI21_X1 port map( B1 => n24, B2 => ENABLE, A => n29, ZN => n19);
   U5 : NAND2_X1 port map( A1 => D(1), A2 => ENABLE, ZN => n29);
   U6 : OAI21_X1 port map( B1 => n23, B2 => ENABLE, A => n28, ZN => n18);
   U7 : NAND2_X1 port map( A1 => D(2), A2 => ENABLE, ZN => n28);
   U8 : OAI21_X1 port map( B1 => n22, B2 => ENABLE, A => n27, ZN => n17);
   U9 : NAND2_X1 port map( A1 => D(3), A2 => ENABLE, ZN => n27);
   U10 : OAI21_X1 port map( B1 => n21, B2 => ENABLE, A => n26, ZN => n16);
   U11 : NAND2_X1 port map( A1 => D(4), A2 => ENABLE, ZN => n26);

end SYN_ASYNCHBEHAV;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FF_7 is

   port( CLK, RESET, EN, D : in std_logic;  Q : out std_logic);

end FF_7;

architecture SYN_SYNC_BHV of FF_7 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n5, n6, n_1034 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFF_X1 port map( D => n5, CK => CLK, Q => Q_port, QN => n_1034);
   U3 : NOR2_X1 port map( A1 => n6, A2 => n1, ZN => n5);
   U4 : AOI22_X1 port map( A1 => EN, A2 => D, B1 => Q_port, B2 => n2, ZN => n6)
                           ;
   U5 : INV_X1 port map( A => EN, ZN => n2);
   U6 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_SYNC_BHV;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FF_6 is

   port( CLK, RESET, EN, D : in std_logic;  Q : out std_logic);

end FF_6;

architecture SYN_SYNC_BHV of FF_6 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n5, n6, n_1035 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFF_X1 port map( D => n5, CK => CLK, Q => Q_port, QN => n_1035);
   U3 : NOR2_X1 port map( A1 => n6, A2 => n1, ZN => n5);
   U4 : AOI22_X1 port map( A1 => EN, A2 => D, B1 => Q_port, B2 => n2, ZN => n6)
                           ;
   U5 : INV_X1 port map( A => EN, ZN => n2);
   U6 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_SYNC_BHV;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FF_5 is

   port( CLK, RESET, EN, D : in std_logic;  Q : out std_logic);

end FF_5;

architecture SYN_SYNC_BHV of FF_5 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n5, n6, n_1036 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFF_X1 port map( D => n5, CK => CLK, Q => Q_port, QN => n_1036);
   U3 : NOR2_X1 port map( A1 => n6, A2 => n1, ZN => n5);
   U4 : AOI22_X1 port map( A1 => EN, A2 => D, B1 => Q_port, B2 => n2, ZN => n6)
                           ;
   U5 : INV_X1 port map( A => EN, ZN => n2);
   U6 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_SYNC_BHV;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FF_4 is

   port( CLK, RESET, EN, D : in std_logic;  Q : out std_logic);

end FF_4;

architecture SYN_SYNC_BHV of FF_4 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component SDFF_X1
      port( D, SI, SE, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n4, n_1037 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : SDFF_X1 port map( D => RESET, SI => n1, SE => n4, CK => CLK, Q => 
                           Q_port, QN => n_1037);
   n1 <= '0';
   U4 : AOI22_X1 port map( A1 => EN, A2 => D, B1 => Q_port, B2 => n2, ZN => n4)
                           ;
   U5 : INV_X1 port map( A => EN, ZN => n2);

end SYN_SYNC_BHV;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FF_3 is

   port( CLK, RESET, EN, D : in std_logic;  Q : out std_logic);

end FF_3;

architecture SYN_SYNC_BHV of FF_3 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n5, n6, n_1038 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFF_X1 port map( D => n5, CK => CLK, Q => Q_port, QN => n_1038);
   U3 : NOR2_X1 port map( A1 => n6, A2 => n1, ZN => n5);
   U4 : AOI22_X1 port map( A1 => EN, A2 => D, B1 => Q_port, B2 => n2, ZN => n6)
                           ;
   U5 : INV_X1 port map( A => EN, ZN => n2);
   U6 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_SYNC_BHV;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FF_2 is

   port( CLK, RESET, EN, D : in std_logic;  Q : out std_logic);

end FF_2;

architecture SYN_SYNC_BHV of FF_2 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n5, n6, n_1039 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFF_X1 port map( D => n5, CK => CLK, Q => Q_port, QN => n_1039);
   U3 : NOR2_X1 port map( A1 => n6, A2 => n1, ZN => n5);
   U4 : AOI22_X1 port map( A1 => EN, A2 => D, B1 => Q_port, B2 => n2, ZN => n6)
                           ;
   U5 : INV_X1 port map( A => EN, ZN => n2);
   U6 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_SYNC_BHV;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FF_1 is

   port( CLK, RESET, EN, D : in std_logic;  Q : out std_logic);

end FF_1;

architecture SYN_SYNC_BHV of FF_1 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n5, n6, n_1040 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFF_X1 port map( D => n5, CK => CLK, Q => Q_port, QN => n_1040);
   U3 : NOR2_X1 port map( A1 => n6, A2 => n1, ZN => n5);
   U4 : AOI22_X1 port map( A1 => EN, A2 => D, B1 => Q_port, B2 => n2, ZN => n6)
                           ;
   U5 : INV_X1 port map( A => EN, ZN => n2);
   U6 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_SYNC_BHV;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_GENERIC_NBIT32_6 is

   port( A, B : in std_logic_vector (31 downto 0);  SEL : in std_logic;  Y : 
         out std_logic_vector (31 downto 0));

end MUX21_GENERIC_NBIT32_6;

architecture SYN_struct of MUX21_GENERIC_NBIT32_6 is

   component MUX21_193
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_194
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_195
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_196
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_197
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_198
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_199
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_200
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_201
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_202
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_203
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_204
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_205
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_206
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_207
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_208
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_209
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_210
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_211
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_212
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_213
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_214
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_215
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_216
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_217
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_218
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_219
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_220
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_221
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_222
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_223
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_224
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;

begin
   
   gen1_0 : MUX21_224 port map( A => A(0), B => B(0), S => SEL, Y => Y(0));
   gen1_1 : MUX21_223 port map( A => A(1), B => B(1), S => SEL, Y => Y(1));
   gen1_2 : MUX21_222 port map( A => A(2), B => B(2), S => SEL, Y => Y(2));
   gen1_3 : MUX21_221 port map( A => A(3), B => B(3), S => SEL, Y => Y(3));
   gen1_4 : MUX21_220 port map( A => A(4), B => B(4), S => SEL, Y => Y(4));
   gen1_5 : MUX21_219 port map( A => A(5), B => B(5), S => SEL, Y => Y(5));
   gen1_6 : MUX21_218 port map( A => A(6), B => B(6), S => SEL, Y => Y(6));
   gen1_7 : MUX21_217 port map( A => A(7), B => B(7), S => SEL, Y => Y(7));
   gen1_8 : MUX21_216 port map( A => A(8), B => B(8), S => SEL, Y => Y(8));
   gen1_9 : MUX21_215 port map( A => A(9), B => B(9), S => SEL, Y => Y(9));
   gen1_10 : MUX21_214 port map( A => A(10), B => B(10), S => SEL, Y => Y(10));
   gen1_11 : MUX21_213 port map( A => A(11), B => B(11), S => SEL, Y => Y(11));
   gen1_12 : MUX21_212 port map( A => A(12), B => B(12), S => SEL, Y => Y(12));
   gen1_13 : MUX21_211 port map( A => A(13), B => B(13), S => SEL, Y => Y(13));
   gen1_14 : MUX21_210 port map( A => A(14), B => B(14), S => SEL, Y => Y(14));
   gen1_15 : MUX21_209 port map( A => A(15), B => B(15), S => SEL, Y => Y(15));
   gen1_16 : MUX21_208 port map( A => A(16), B => B(16), S => SEL, Y => Y(16));
   gen1_17 : MUX21_207 port map( A => A(17), B => B(17), S => SEL, Y => Y(17));
   gen1_18 : MUX21_206 port map( A => A(18), B => B(18), S => SEL, Y => Y(18));
   gen1_19 : MUX21_205 port map( A => A(19), B => B(19), S => SEL, Y => Y(19));
   gen1_20 : MUX21_204 port map( A => A(20), B => B(20), S => SEL, Y => Y(20));
   gen1_21 : MUX21_203 port map( A => A(21), B => B(21), S => SEL, Y => Y(21));
   gen1_22 : MUX21_202 port map( A => A(22), B => B(22), S => SEL, Y => Y(22));
   gen1_23 : MUX21_201 port map( A => A(23), B => B(23), S => SEL, Y => Y(23));
   gen1_24 : MUX21_200 port map( A => A(24), B => B(24), S => SEL, Y => Y(24));
   gen1_25 : MUX21_199 port map( A => A(25), B => B(25), S => SEL, Y => Y(25));
   gen1_26 : MUX21_198 port map( A => A(26), B => B(26), S => SEL, Y => Y(26));
   gen1_27 : MUX21_197 port map( A => A(27), B => B(27), S => SEL, Y => Y(27));
   gen1_28 : MUX21_196 port map( A => A(28), B => B(28), S => SEL, Y => Y(28));
   gen1_29 : MUX21_195 port map( A => A(29), B => B(29), S => SEL, Y => Y(29));
   gen1_30 : MUX21_194 port map( A => A(30), B => B(30), S => SEL, Y => Y(30));
   gen1_31 : MUX21_193 port map( A => A(31), B => B(31), S => SEL, Y => Y(31));

end SYN_struct;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_GENERIC_NBIT32_5 is

   port( A, B : in std_logic_vector (31 downto 0);  SEL : in std_logic;  Y : 
         out std_logic_vector (31 downto 0));

end MUX21_GENERIC_NBIT32_5;

architecture SYN_struct of MUX21_GENERIC_NBIT32_5 is

   component MUX21_161
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_162
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_163
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_164
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_165
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_166
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_167
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_168
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_169
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_170
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_171
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_172
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_173
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_174
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_175
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_176
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_177
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_178
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_179
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_180
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_181
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_182
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_183
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_184
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_185
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_186
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_187
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_188
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_189
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_190
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_191
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_192
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;

begin
   
   gen1_0 : MUX21_192 port map( A => A(0), B => B(0), S => SEL, Y => Y(0));
   gen1_1 : MUX21_191 port map( A => A(1), B => B(1), S => SEL, Y => Y(1));
   gen1_2 : MUX21_190 port map( A => A(2), B => B(2), S => SEL, Y => Y(2));
   gen1_3 : MUX21_189 port map( A => A(3), B => B(3), S => SEL, Y => Y(3));
   gen1_4 : MUX21_188 port map( A => A(4), B => B(4), S => SEL, Y => Y(4));
   gen1_5 : MUX21_187 port map( A => A(5), B => B(5), S => SEL, Y => Y(5));
   gen1_6 : MUX21_186 port map( A => A(6), B => B(6), S => SEL, Y => Y(6));
   gen1_7 : MUX21_185 port map( A => A(7), B => B(7), S => SEL, Y => Y(7));
   gen1_8 : MUX21_184 port map( A => A(8), B => B(8), S => SEL, Y => Y(8));
   gen1_9 : MUX21_183 port map( A => A(9), B => B(9), S => SEL, Y => Y(9));
   gen1_10 : MUX21_182 port map( A => A(10), B => B(10), S => SEL, Y => Y(10));
   gen1_11 : MUX21_181 port map( A => A(11), B => B(11), S => SEL, Y => Y(11));
   gen1_12 : MUX21_180 port map( A => A(12), B => B(12), S => SEL, Y => Y(12));
   gen1_13 : MUX21_179 port map( A => A(13), B => B(13), S => SEL, Y => Y(13));
   gen1_14 : MUX21_178 port map( A => A(14), B => B(14), S => SEL, Y => Y(14));
   gen1_15 : MUX21_177 port map( A => A(15), B => B(15), S => SEL, Y => Y(15));
   gen1_16 : MUX21_176 port map( A => A(16), B => B(16), S => SEL, Y => Y(16));
   gen1_17 : MUX21_175 port map( A => A(17), B => B(17), S => SEL, Y => Y(17));
   gen1_18 : MUX21_174 port map( A => A(18), B => B(18), S => SEL, Y => Y(18));
   gen1_19 : MUX21_173 port map( A => A(19), B => B(19), S => SEL, Y => Y(19));
   gen1_20 : MUX21_172 port map( A => A(20), B => B(20), S => SEL, Y => Y(20));
   gen1_21 : MUX21_171 port map( A => A(21), B => B(21), S => SEL, Y => Y(21));
   gen1_22 : MUX21_170 port map( A => A(22), B => B(22), S => SEL, Y => Y(22));
   gen1_23 : MUX21_169 port map( A => A(23), B => B(23), S => SEL, Y => Y(23));
   gen1_24 : MUX21_168 port map( A => A(24), B => B(24), S => SEL, Y => Y(24));
   gen1_25 : MUX21_167 port map( A => A(25), B => B(25), S => SEL, Y => Y(25));
   gen1_26 : MUX21_166 port map( A => A(26), B => B(26), S => SEL, Y => Y(26));
   gen1_27 : MUX21_165 port map( A => A(27), B => B(27), S => SEL, Y => Y(27));
   gen1_28 : MUX21_164 port map( A => A(28), B => B(28), S => SEL, Y => Y(28));
   gen1_29 : MUX21_163 port map( A => A(29), B => B(29), S => SEL, Y => Y(29));
   gen1_30 : MUX21_162 port map( A => A(30), B => B(30), S => SEL, Y => Y(30));
   gen1_31 : MUX21_161 port map( A => A(31), B => B(31), S => SEL, Y => Y(31));

end SYN_struct;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_GENERIC_NBIT32_4 is

   port( A, B : in std_logic_vector (31 downto 0);  SEL : in std_logic;  Y : 
         out std_logic_vector (31 downto 0));

end MUX21_GENERIC_NBIT32_4;

architecture SYN_struct of MUX21_GENERIC_NBIT32_4 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component MUX21_129
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_130
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_131
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_132
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_133
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_134
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_135
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_136
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_137
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_138
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_139
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_140
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_141
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_142
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_143
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_144
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_145
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_146
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_147
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_148
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_149
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_150
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_151
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_152
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_153
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_154
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_155
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_156
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_157
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_158
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_159
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_160
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   signal n1, n2, n3 : std_logic;

begin
   
   gen1_0 : MUX21_160 port map( A => A(0), B => B(0), S => n1, Y => Y(0));
   gen1_1 : MUX21_159 port map( A => A(1), B => B(1), S => n1, Y => Y(1));
   gen1_2 : MUX21_158 port map( A => A(2), B => B(2), S => n1, Y => Y(2));
   gen1_3 : MUX21_157 port map( A => A(3), B => B(3), S => n1, Y => Y(3));
   gen1_4 : MUX21_156 port map( A => A(4), B => B(4), S => n1, Y => Y(4));
   gen1_5 : MUX21_155 port map( A => A(5), B => B(5), S => n1, Y => Y(5));
   gen1_6 : MUX21_154 port map( A => A(6), B => B(6), S => n1, Y => Y(6));
   gen1_7 : MUX21_153 port map( A => A(7), B => B(7), S => n1, Y => Y(7));
   gen1_8 : MUX21_152 port map( A => A(8), B => B(8), S => n1, Y => Y(8));
   gen1_9 : MUX21_151 port map( A => A(9), B => B(9), S => n1, Y => Y(9));
   gen1_10 : MUX21_150 port map( A => A(10), B => B(10), S => n1, Y => Y(10));
   gen1_11 : MUX21_149 port map( A => A(11), B => B(11), S => n1, Y => Y(11));
   gen1_12 : MUX21_148 port map( A => A(12), B => B(12), S => n2, Y => Y(12));
   gen1_13 : MUX21_147 port map( A => A(13), B => B(13), S => n2, Y => Y(13));
   gen1_14 : MUX21_146 port map( A => A(14), B => B(14), S => n2, Y => Y(14));
   gen1_15 : MUX21_145 port map( A => A(15), B => B(15), S => n2, Y => Y(15));
   gen1_16 : MUX21_144 port map( A => A(16), B => B(16), S => n2, Y => Y(16));
   gen1_17 : MUX21_143 port map( A => A(17), B => B(17), S => n2, Y => Y(17));
   gen1_18 : MUX21_142 port map( A => A(18), B => B(18), S => n2, Y => Y(18));
   gen1_19 : MUX21_141 port map( A => A(19), B => B(19), S => n2, Y => Y(19));
   gen1_20 : MUX21_140 port map( A => A(20), B => B(20), S => n2, Y => Y(20));
   gen1_21 : MUX21_139 port map( A => A(21), B => B(21), S => n2, Y => Y(21));
   gen1_22 : MUX21_138 port map( A => A(22), B => B(22), S => n2, Y => Y(22));
   gen1_23 : MUX21_137 port map( A => A(23), B => B(23), S => n2, Y => Y(23));
   gen1_24 : MUX21_136 port map( A => A(24), B => B(24), S => n3, Y => Y(24));
   gen1_25 : MUX21_135 port map( A => A(25), B => B(25), S => n3, Y => Y(25));
   gen1_26 : MUX21_134 port map( A => A(26), B => B(26), S => n3, Y => Y(26));
   gen1_27 : MUX21_133 port map( A => A(27), B => B(27), S => n3, Y => Y(27));
   gen1_28 : MUX21_132 port map( A => A(28), B => B(28), S => n3, Y => Y(28));
   gen1_29 : MUX21_131 port map( A => A(29), B => B(29), S => n3, Y => Y(29));
   gen1_30 : MUX21_130 port map( A => A(30), B => B(30), S => n3, Y => Y(30));
   gen1_31 : MUX21_129 port map( A => A(31), B => B(31), S => n3, Y => Y(31));
   U1 : BUF_X1 port map( A => SEL, Z => n1);
   U2 : BUF_X1 port map( A => SEL, Z => n2);
   U3 : BUF_X1 port map( A => SEL, Z => n3);

end SYN_struct;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_GENERIC_NBIT32_3 is

   port( A, B : in std_logic_vector (31 downto 0);  SEL : in std_logic;  Y : 
         out std_logic_vector (31 downto 0));

end MUX21_GENERIC_NBIT32_3;

architecture SYN_struct of MUX21_GENERIC_NBIT32_3 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component MUX21_97
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_98
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_99
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_100
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_101
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_102
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_103
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_104
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_105
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_106
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_107
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_108
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_109
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_110
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_111
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_112
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_113
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_114
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_115
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_116
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_117
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_118
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_119
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_120
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_121
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_122
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_123
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_124
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_125
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_126
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_127
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_128
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   signal n1, n2, n3 : std_logic;

begin
   
   gen1_0 : MUX21_128 port map( A => A(0), B => B(0), S => n1, Y => Y(0));
   gen1_1 : MUX21_127 port map( A => A(1), B => B(1), S => n1, Y => Y(1));
   gen1_2 : MUX21_126 port map( A => A(2), B => B(2), S => n1, Y => Y(2));
   gen1_3 : MUX21_125 port map( A => A(3), B => B(3), S => n1, Y => Y(3));
   gen1_4 : MUX21_124 port map( A => A(4), B => B(4), S => n1, Y => Y(4));
   gen1_5 : MUX21_123 port map( A => A(5), B => B(5), S => n1, Y => Y(5));
   gen1_6 : MUX21_122 port map( A => A(6), B => B(6), S => n1, Y => Y(6));
   gen1_7 : MUX21_121 port map( A => A(7), B => B(7), S => n1, Y => Y(7));
   gen1_8 : MUX21_120 port map( A => A(8), B => B(8), S => n1, Y => Y(8));
   gen1_9 : MUX21_119 port map( A => A(9), B => B(9), S => n1, Y => Y(9));
   gen1_10 : MUX21_118 port map( A => A(10), B => B(10), S => n1, Y => Y(10));
   gen1_11 : MUX21_117 port map( A => A(11), B => B(11), S => n1, Y => Y(11));
   gen1_12 : MUX21_116 port map( A => A(12), B => B(12), S => n2, Y => Y(12));
   gen1_13 : MUX21_115 port map( A => A(13), B => B(13), S => n2, Y => Y(13));
   gen1_14 : MUX21_114 port map( A => A(14), B => B(14), S => n2, Y => Y(14));
   gen1_15 : MUX21_113 port map( A => A(15), B => B(15), S => n2, Y => Y(15));
   gen1_16 : MUX21_112 port map( A => A(16), B => B(16), S => n2, Y => Y(16));
   gen1_17 : MUX21_111 port map( A => A(17), B => B(17), S => n2, Y => Y(17));
   gen1_18 : MUX21_110 port map( A => A(18), B => B(18), S => n2, Y => Y(18));
   gen1_19 : MUX21_109 port map( A => A(19), B => B(19), S => n2, Y => Y(19));
   gen1_20 : MUX21_108 port map( A => A(20), B => B(20), S => n2, Y => Y(20));
   gen1_21 : MUX21_107 port map( A => A(21), B => B(21), S => n2, Y => Y(21));
   gen1_22 : MUX21_106 port map( A => A(22), B => B(22), S => n2, Y => Y(22));
   gen1_23 : MUX21_105 port map( A => A(23), B => B(23), S => n2, Y => Y(23));
   gen1_24 : MUX21_104 port map( A => A(24), B => B(24), S => n3, Y => Y(24));
   gen1_25 : MUX21_103 port map( A => A(25), B => B(25), S => n3, Y => Y(25));
   gen1_26 : MUX21_102 port map( A => A(26), B => B(26), S => n3, Y => Y(26));
   gen1_27 : MUX21_101 port map( A => A(27), B => B(27), S => n3, Y => Y(27));
   gen1_28 : MUX21_100 port map( A => A(28), B => B(28), S => n3, Y => Y(28));
   gen1_29 : MUX21_99 port map( A => A(29), B => B(29), S => n3, Y => Y(29));
   gen1_30 : MUX21_98 port map( A => A(30), B => B(30), S => n3, Y => Y(30));
   gen1_31 : MUX21_97 port map( A => A(31), B => B(31), S => n3, Y => Y(31));
   U1 : BUF_X1 port map( A => SEL, Z => n1);
   U2 : BUF_X1 port map( A => SEL, Z => n2);
   U3 : BUF_X1 port map( A => SEL, Z => n3);

end SYN_struct;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_GENERIC_NBIT32_2 is

   port( A, B : in std_logic_vector (31 downto 0);  SEL : in std_logic;  Y : 
         out std_logic_vector (31 downto 0));

end MUX21_GENERIC_NBIT32_2;

architecture SYN_struct of MUX21_GENERIC_NBIT32_2 is

   component MUX21_65
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_66
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_67
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_68
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_69
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_70
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_71
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_72
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_73
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_74
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_75
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_76
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_77
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_78
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_79
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_80
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_81
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_82
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_83
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_84
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_85
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_86
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_87
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_88
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_89
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_90
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_91
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_92
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_93
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_94
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_95
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_96
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;

begin
   
   gen1_0 : MUX21_96 port map( A => A(0), B => B(0), S => SEL, Y => Y(0));
   gen1_1 : MUX21_95 port map( A => A(1), B => B(1), S => SEL, Y => Y(1));
   gen1_2 : MUX21_94 port map( A => A(2), B => B(2), S => SEL, Y => Y(2));
   gen1_3 : MUX21_93 port map( A => A(3), B => B(3), S => SEL, Y => Y(3));
   gen1_4 : MUX21_92 port map( A => A(4), B => B(4), S => SEL, Y => Y(4));
   gen1_5 : MUX21_91 port map( A => A(5), B => B(5), S => SEL, Y => Y(5));
   gen1_6 : MUX21_90 port map( A => A(6), B => B(6), S => SEL, Y => Y(6));
   gen1_7 : MUX21_89 port map( A => A(7), B => B(7), S => SEL, Y => Y(7));
   gen1_8 : MUX21_88 port map( A => A(8), B => B(8), S => SEL, Y => Y(8));
   gen1_9 : MUX21_87 port map( A => A(9), B => B(9), S => SEL, Y => Y(9));
   gen1_10 : MUX21_86 port map( A => A(10), B => B(10), S => SEL, Y => Y(10));
   gen1_11 : MUX21_85 port map( A => A(11), B => B(11), S => SEL, Y => Y(11));
   gen1_12 : MUX21_84 port map( A => A(12), B => B(12), S => SEL, Y => Y(12));
   gen1_13 : MUX21_83 port map( A => A(13), B => B(13), S => SEL, Y => Y(13));
   gen1_14 : MUX21_82 port map( A => A(14), B => B(14), S => SEL, Y => Y(14));
   gen1_15 : MUX21_81 port map( A => A(15), B => B(15), S => SEL, Y => Y(15));
   gen1_16 : MUX21_80 port map( A => A(16), B => B(16), S => SEL, Y => Y(16));
   gen1_17 : MUX21_79 port map( A => A(17), B => B(17), S => SEL, Y => Y(17));
   gen1_18 : MUX21_78 port map( A => A(18), B => B(18), S => SEL, Y => Y(18));
   gen1_19 : MUX21_77 port map( A => A(19), B => B(19), S => SEL, Y => Y(19));
   gen1_20 : MUX21_76 port map( A => A(20), B => B(20), S => SEL, Y => Y(20));
   gen1_21 : MUX21_75 port map( A => A(21), B => B(21), S => SEL, Y => Y(21));
   gen1_22 : MUX21_74 port map( A => A(22), B => B(22), S => SEL, Y => Y(22));
   gen1_23 : MUX21_73 port map( A => A(23), B => B(23), S => SEL, Y => Y(23));
   gen1_24 : MUX21_72 port map( A => A(24), B => B(24), S => SEL, Y => Y(24));
   gen1_25 : MUX21_71 port map( A => A(25), B => B(25), S => SEL, Y => Y(25));
   gen1_26 : MUX21_70 port map( A => A(26), B => B(26), S => SEL, Y => Y(26));
   gen1_27 : MUX21_69 port map( A => A(27), B => B(27), S => SEL, Y => Y(27));
   gen1_28 : MUX21_68 port map( A => A(28), B => B(28), S => SEL, Y => Y(28));
   gen1_29 : MUX21_67 port map( A => A(29), B => B(29), S => SEL, Y => Y(29));
   gen1_30 : MUX21_66 port map( A => A(30), B => B(30), S => SEL, Y => Y(30));
   gen1_31 : MUX21_65 port map( A => A(31), B => B(31), S => SEL, Y => Y(31));

end SYN_struct;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_GENERIC_NBIT32_1 is

   port( A, B : in std_logic_vector (31 downto 0);  SEL : in std_logic;  Y : 
         out std_logic_vector (31 downto 0));

end MUX21_GENERIC_NBIT32_1;

architecture SYN_struct of MUX21_GENERIC_NBIT32_1 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component MUX21_33
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_34
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_35
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_36
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_37
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_38
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_39
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_40
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_41
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_42
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_43
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_44
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_45
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_46
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_47
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_48
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_49
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_50
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_51
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_52
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_53
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_54
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_55
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_56
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_57
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_58
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_59
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_60
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_61
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_62
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_63
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_64
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   signal n1, n2, n3 : std_logic;

begin
   
   gen1_0 : MUX21_64 port map( A => A(0), B => B(0), S => n1, Y => Y(0));
   gen1_1 : MUX21_63 port map( A => A(1), B => B(1), S => n1, Y => Y(1));
   gen1_2 : MUX21_62 port map( A => A(2), B => B(2), S => n1, Y => Y(2));
   gen1_3 : MUX21_61 port map( A => A(3), B => B(3), S => n1, Y => Y(3));
   gen1_4 : MUX21_60 port map( A => A(4), B => B(4), S => n1, Y => Y(4));
   gen1_5 : MUX21_59 port map( A => A(5), B => B(5), S => n1, Y => Y(5));
   gen1_6 : MUX21_58 port map( A => A(6), B => B(6), S => n1, Y => Y(6));
   gen1_7 : MUX21_57 port map( A => A(7), B => B(7), S => n1, Y => Y(7));
   gen1_8 : MUX21_56 port map( A => A(8), B => B(8), S => n1, Y => Y(8));
   gen1_9 : MUX21_55 port map( A => A(9), B => B(9), S => n1, Y => Y(9));
   gen1_10 : MUX21_54 port map( A => A(10), B => B(10), S => n1, Y => Y(10));
   gen1_11 : MUX21_53 port map( A => A(11), B => B(11), S => n1, Y => Y(11));
   gen1_12 : MUX21_52 port map( A => A(12), B => B(12), S => n2, Y => Y(12));
   gen1_13 : MUX21_51 port map( A => A(13), B => B(13), S => n2, Y => Y(13));
   gen1_14 : MUX21_50 port map( A => A(14), B => B(14), S => n2, Y => Y(14));
   gen1_15 : MUX21_49 port map( A => A(15), B => B(15), S => n2, Y => Y(15));
   gen1_16 : MUX21_48 port map( A => A(16), B => B(16), S => n2, Y => Y(16));
   gen1_17 : MUX21_47 port map( A => A(17), B => B(17), S => n2, Y => Y(17));
   gen1_18 : MUX21_46 port map( A => A(18), B => B(18), S => n2, Y => Y(18));
   gen1_19 : MUX21_45 port map( A => A(19), B => B(19), S => n2, Y => Y(19));
   gen1_20 : MUX21_44 port map( A => A(20), B => B(20), S => n2, Y => Y(20));
   gen1_21 : MUX21_43 port map( A => A(21), B => B(21), S => n2, Y => Y(21));
   gen1_22 : MUX21_42 port map( A => A(22), B => B(22), S => n2, Y => Y(22));
   gen1_23 : MUX21_41 port map( A => A(23), B => B(23), S => n2, Y => Y(23));
   gen1_24 : MUX21_40 port map( A => A(24), B => B(24), S => n3, Y => Y(24));
   gen1_25 : MUX21_39 port map( A => A(25), B => B(25), S => n3, Y => Y(25));
   gen1_26 : MUX21_38 port map( A => A(26), B => B(26), S => n3, Y => Y(26));
   gen1_27 : MUX21_37 port map( A => A(27), B => B(27), S => n3, Y => Y(27));
   gen1_28 : MUX21_36 port map( A => A(28), B => B(28), S => n3, Y => Y(28));
   gen1_29 : MUX21_35 port map( A => A(29), B => B(29), S => n3, Y => Y(29));
   gen1_30 : MUX21_34 port map( A => A(30), B => B(30), S => n3, Y => Y(30));
   gen1_31 : MUX21_33 port map( A => A(31), B => B(31), S => n3, Y => Y(31));
   U1 : BUF_X1 port map( A => SEL, Z => n1);
   U2 : BUF_X1 port map( A => SEL, Z => n2);
   U3 : BUF_X1 port map( A => SEL, Z => n3);

end SYN_struct;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity regFFD_NBIT32_18 is

   port( CK, RESET, ENABLE : in std_logic;  D : in std_logic_vector (31 downto 
         0);  Q : out std_logic_vector (31 downto 0));

end regFFD_NBIT32_18;

architecture SYN_ASYNCHBEHAV of regFFD_NBIT32_18 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, 
      n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, 
      n121, n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, 
      n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, 
      n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, 
      n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, 
      n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, 
      n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, 
      n193, n194, n195 : std_logic;

begin
   
   Q_reg_31_inst : DFFR_X1 port map( D => n100, CK => CK, RN => n99, Q => Q(31)
                           , QN => n132);
   Q_reg_30_inst : DFFR_X1 port map( D => n101, CK => CK, RN => n99, Q => Q(30)
                           , QN => n133);
   Q_reg_29_inst : DFFR_X1 port map( D => n102, CK => CK, RN => n99, Q => Q(29)
                           , QN => n134);
   Q_reg_28_inst : DFFR_X1 port map( D => n103, CK => CK, RN => n99, Q => Q(28)
                           , QN => n135);
   Q_reg_27_inst : DFFR_X1 port map( D => n104, CK => CK, RN => n99, Q => Q(27)
                           , QN => n136);
   Q_reg_26_inst : DFFR_X1 port map( D => n105, CK => CK, RN => n99, Q => Q(26)
                           , QN => n137);
   Q_reg_25_inst : DFFR_X1 port map( D => n106, CK => CK, RN => n99, Q => Q(25)
                           , QN => n138);
   Q_reg_24_inst : DFFR_X1 port map( D => n107, CK => CK, RN => n99, Q => Q(24)
                           , QN => n139);
   Q_reg_23_inst : DFFR_X1 port map( D => n108, CK => CK, RN => n98, Q => Q(23)
                           , QN => n140);
   Q_reg_22_inst : DFFR_X1 port map( D => n109, CK => CK, RN => n98, Q => Q(22)
                           , QN => n141);
   Q_reg_21_inst : DFFR_X1 port map( D => n110, CK => CK, RN => n98, Q => Q(21)
                           , QN => n142);
   Q_reg_20_inst : DFFR_X1 port map( D => n111, CK => CK, RN => n98, Q => Q(20)
                           , QN => n143);
   Q_reg_19_inst : DFFR_X1 port map( D => n112, CK => CK, RN => n98, Q => Q(19)
                           , QN => n144);
   Q_reg_18_inst : DFFR_X1 port map( D => n113, CK => CK, RN => n98, Q => Q(18)
                           , QN => n145);
   Q_reg_17_inst : DFFR_X1 port map( D => n114, CK => CK, RN => n98, Q => Q(17)
                           , QN => n146);
   Q_reg_16_inst : DFFR_X1 port map( D => n115, CK => CK, RN => n98, Q => Q(16)
                           , QN => n147);
   Q_reg_15_inst : DFFR_X1 port map( D => n116, CK => CK, RN => n98, Q => Q(15)
                           , QN => n148);
   Q_reg_14_inst : DFFR_X1 port map( D => n117, CK => CK, RN => n98, Q => Q(14)
                           , QN => n149);
   Q_reg_13_inst : DFFR_X1 port map( D => n118, CK => CK, RN => n98, Q => Q(13)
                           , QN => n150);
   Q_reg_12_inst : DFFR_X1 port map( D => n119, CK => CK, RN => n98, Q => Q(12)
                           , QN => n151);
   Q_reg_11_inst : DFFR_X1 port map( D => n120, CK => CK, RN => n97, Q => Q(11)
                           , QN => n152);
   Q_reg_10_inst : DFFR_X1 port map( D => n121, CK => CK, RN => n97, Q => Q(10)
                           , QN => n153);
   Q_reg_9_inst : DFFR_X1 port map( D => n122, CK => CK, RN => n97, Q => Q(9), 
                           QN => n154);
   Q_reg_8_inst : DFFR_X1 port map( D => n123, CK => CK, RN => n97, Q => Q(8), 
                           QN => n155);
   Q_reg_7_inst : DFFR_X1 port map( D => n124, CK => CK, RN => n97, Q => Q(7), 
                           QN => n156);
   Q_reg_6_inst : DFFR_X1 port map( D => n125, CK => CK, RN => n97, Q => Q(6), 
                           QN => n157);
   Q_reg_5_inst : DFFR_X1 port map( D => n126, CK => CK, RN => n97, Q => Q(5), 
                           QN => n158);
   Q_reg_4_inst : DFFR_X1 port map( D => n127, CK => CK, RN => n97, Q => Q(4), 
                           QN => n159);
   Q_reg_3_inst : DFFR_X1 port map( D => n128, CK => CK, RN => n97, Q => Q(3), 
                           QN => n160);
   Q_reg_2_inst : DFFR_X1 port map( D => n129, CK => CK, RN => n97, Q => Q(2), 
                           QN => n161);
   Q_reg_1_inst : DFFR_X1 port map( D => n130, CK => CK, RN => n97, Q => Q(1), 
                           QN => n162);
   Q_reg_0_inst : DFFR_X1 port map( D => n131, CK => CK, RN => n97, Q => Q(0), 
                           QN => n163);
   U2 : BUF_X1 port map( A => RESET, Z => n97);
   U3 : BUF_X1 port map( A => RESET, Z => n98);
   U4 : BUF_X1 port map( A => RESET, Z => n99);
   U5 : OAI21_X1 port map( B1 => n163, B2 => ENABLE, A => n195, ZN => n131);
   U6 : NAND2_X1 port map( A1 => ENABLE, A2 => D(0), ZN => n195);
   U7 : OAI21_X1 port map( B1 => n162, B2 => ENABLE, A => n194, ZN => n130);
   U8 : NAND2_X1 port map( A1 => D(1), A2 => ENABLE, ZN => n194);
   U9 : OAI21_X1 port map( B1 => n161, B2 => ENABLE, A => n193, ZN => n129);
   U10 : NAND2_X1 port map( A1 => D(2), A2 => ENABLE, ZN => n193);
   U11 : OAI21_X1 port map( B1 => n160, B2 => ENABLE, A => n192, ZN => n128);
   U12 : NAND2_X1 port map( A1 => D(3), A2 => ENABLE, ZN => n192);
   U13 : OAI21_X1 port map( B1 => n159, B2 => ENABLE, A => n191, ZN => n127);
   U14 : NAND2_X1 port map( A1 => D(4), A2 => ENABLE, ZN => n191);
   U15 : OAI21_X1 port map( B1 => n158, B2 => ENABLE, A => n190, ZN => n126);
   U16 : NAND2_X1 port map( A1 => D(5), A2 => ENABLE, ZN => n190);
   U17 : OAI21_X1 port map( B1 => n157, B2 => ENABLE, A => n189, ZN => n125);
   U18 : NAND2_X1 port map( A1 => D(6), A2 => ENABLE, ZN => n189);
   U19 : OAI21_X1 port map( B1 => n156, B2 => ENABLE, A => n188, ZN => n124);
   U20 : NAND2_X1 port map( A1 => D(7), A2 => ENABLE, ZN => n188);
   U21 : OAI21_X1 port map( B1 => n155, B2 => ENABLE, A => n187, ZN => n123);
   U22 : NAND2_X1 port map( A1 => D(8), A2 => ENABLE, ZN => n187);
   U23 : OAI21_X1 port map( B1 => n154, B2 => ENABLE, A => n186, ZN => n122);
   U24 : NAND2_X1 port map( A1 => D(9), A2 => ENABLE, ZN => n186);
   U25 : OAI21_X1 port map( B1 => n153, B2 => ENABLE, A => n185, ZN => n121);
   U26 : NAND2_X1 port map( A1 => D(10), A2 => ENABLE, ZN => n185);
   U27 : OAI21_X1 port map( B1 => n152, B2 => ENABLE, A => n184, ZN => n120);
   U28 : NAND2_X1 port map( A1 => D(11), A2 => ENABLE, ZN => n184);
   U29 : OAI21_X1 port map( B1 => n151, B2 => ENABLE, A => n183, ZN => n119);
   U30 : NAND2_X1 port map( A1 => D(12), A2 => ENABLE, ZN => n183);
   U31 : OAI21_X1 port map( B1 => n150, B2 => ENABLE, A => n182, ZN => n118);
   U32 : NAND2_X1 port map( A1 => D(13), A2 => ENABLE, ZN => n182);
   U33 : OAI21_X1 port map( B1 => n149, B2 => ENABLE, A => n181, ZN => n117);
   U34 : NAND2_X1 port map( A1 => D(14), A2 => ENABLE, ZN => n181);
   U35 : OAI21_X1 port map( B1 => n148, B2 => ENABLE, A => n180, ZN => n116);
   U36 : NAND2_X1 port map( A1 => D(15), A2 => ENABLE, ZN => n180);
   U37 : OAI21_X1 port map( B1 => n147, B2 => ENABLE, A => n179, ZN => n115);
   U38 : NAND2_X1 port map( A1 => D(16), A2 => ENABLE, ZN => n179);
   U39 : OAI21_X1 port map( B1 => n146, B2 => ENABLE, A => n178, ZN => n114);
   U40 : NAND2_X1 port map( A1 => D(17), A2 => ENABLE, ZN => n178);
   U41 : OAI21_X1 port map( B1 => n145, B2 => ENABLE, A => n177, ZN => n113);
   U42 : NAND2_X1 port map( A1 => D(18), A2 => ENABLE, ZN => n177);
   U43 : OAI21_X1 port map( B1 => n144, B2 => ENABLE, A => n176, ZN => n112);
   U44 : NAND2_X1 port map( A1 => D(19), A2 => ENABLE, ZN => n176);
   U45 : OAI21_X1 port map( B1 => n143, B2 => ENABLE, A => n175, ZN => n111);
   U46 : NAND2_X1 port map( A1 => D(20), A2 => ENABLE, ZN => n175);
   U47 : OAI21_X1 port map( B1 => n142, B2 => ENABLE, A => n174, ZN => n110);
   U48 : NAND2_X1 port map( A1 => D(21), A2 => ENABLE, ZN => n174);
   U49 : OAI21_X1 port map( B1 => n141, B2 => ENABLE, A => n173, ZN => n109);
   U50 : NAND2_X1 port map( A1 => D(22), A2 => ENABLE, ZN => n173);
   U51 : OAI21_X1 port map( B1 => n140, B2 => ENABLE, A => n172, ZN => n108);
   U52 : NAND2_X1 port map( A1 => D(23), A2 => ENABLE, ZN => n172);
   U53 : OAI21_X1 port map( B1 => n139, B2 => ENABLE, A => n171, ZN => n107);
   U54 : NAND2_X1 port map( A1 => D(24), A2 => ENABLE, ZN => n171);
   U55 : OAI21_X1 port map( B1 => n138, B2 => ENABLE, A => n170, ZN => n106);
   U56 : NAND2_X1 port map( A1 => D(25), A2 => ENABLE, ZN => n170);
   U57 : OAI21_X1 port map( B1 => n137, B2 => ENABLE, A => n169, ZN => n105);
   U58 : NAND2_X1 port map( A1 => D(26), A2 => ENABLE, ZN => n169);
   U59 : OAI21_X1 port map( B1 => n136, B2 => ENABLE, A => n168, ZN => n104);
   U60 : NAND2_X1 port map( A1 => D(27), A2 => ENABLE, ZN => n168);
   U61 : OAI21_X1 port map( B1 => n135, B2 => ENABLE, A => n167, ZN => n103);
   U62 : NAND2_X1 port map( A1 => D(28), A2 => ENABLE, ZN => n167);
   U63 : OAI21_X1 port map( B1 => n134, B2 => ENABLE, A => n166, ZN => n102);
   U64 : NAND2_X1 port map( A1 => D(29), A2 => ENABLE, ZN => n166);
   U65 : OAI21_X1 port map( B1 => n133, B2 => ENABLE, A => n165, ZN => n101);
   U66 : NAND2_X1 port map( A1 => D(30), A2 => ENABLE, ZN => n165);
   U67 : OAI21_X1 port map( B1 => n132, B2 => ENABLE, A => n164, ZN => n100);
   U68 : NAND2_X1 port map( A1 => D(31), A2 => ENABLE, ZN => n164);

end SYN_ASYNCHBEHAV;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity regFFD_NBIT32_17 is

   port( CK, RESET, ENABLE : in std_logic;  D : in std_logic_vector (31 downto 
         0);  Q : out std_logic_vector (31 downto 0));

end regFFD_NBIT32_17;

architecture SYN_ASYNCHBEHAV of regFFD_NBIT32_17 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, 
      n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, 
      n121, n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, 
      n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, 
      n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, 
      n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, 
      n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, 
      n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, 
      n193, n194, n195 : std_logic;

begin
   
   Q_reg_31_inst : DFFR_X1 port map( D => n100, CK => CK, RN => n99, Q => Q(31)
                           , QN => n132);
   Q_reg_30_inst : DFFR_X1 port map( D => n101, CK => CK, RN => n99, Q => Q(30)
                           , QN => n133);
   Q_reg_29_inst : DFFR_X1 port map( D => n102, CK => CK, RN => n99, Q => Q(29)
                           , QN => n134);
   Q_reg_28_inst : DFFR_X1 port map( D => n103, CK => CK, RN => n99, Q => Q(28)
                           , QN => n135);
   Q_reg_27_inst : DFFR_X1 port map( D => n104, CK => CK, RN => n99, Q => Q(27)
                           , QN => n136);
   Q_reg_26_inst : DFFR_X1 port map( D => n105, CK => CK, RN => n99, Q => Q(26)
                           , QN => n137);
   Q_reg_25_inst : DFFR_X1 port map( D => n106, CK => CK, RN => n99, Q => Q(25)
                           , QN => n138);
   Q_reg_24_inst : DFFR_X1 port map( D => n107, CK => CK, RN => n99, Q => Q(24)
                           , QN => n139);
   Q_reg_23_inst : DFFR_X1 port map( D => n108, CK => CK, RN => n98, Q => Q(23)
                           , QN => n140);
   Q_reg_22_inst : DFFR_X1 port map( D => n109, CK => CK, RN => n98, Q => Q(22)
                           , QN => n141);
   Q_reg_21_inst : DFFR_X1 port map( D => n110, CK => CK, RN => n98, Q => Q(21)
                           , QN => n142);
   Q_reg_20_inst : DFFR_X1 port map( D => n111, CK => CK, RN => n98, Q => Q(20)
                           , QN => n143);
   Q_reg_19_inst : DFFR_X1 port map( D => n112, CK => CK, RN => n98, Q => Q(19)
                           , QN => n144);
   Q_reg_18_inst : DFFR_X1 port map( D => n113, CK => CK, RN => n98, Q => Q(18)
                           , QN => n145);
   Q_reg_17_inst : DFFR_X1 port map( D => n114, CK => CK, RN => n98, Q => Q(17)
                           , QN => n146);
   Q_reg_16_inst : DFFR_X1 port map( D => n115, CK => CK, RN => n98, Q => Q(16)
                           , QN => n147);
   Q_reg_15_inst : DFFR_X1 port map( D => n116, CK => CK, RN => n98, Q => Q(15)
                           , QN => n148);
   Q_reg_14_inst : DFFR_X1 port map( D => n117, CK => CK, RN => n98, Q => Q(14)
                           , QN => n149);
   Q_reg_13_inst : DFFR_X1 port map( D => n118, CK => CK, RN => n98, Q => Q(13)
                           , QN => n150);
   Q_reg_12_inst : DFFR_X1 port map( D => n119, CK => CK, RN => n98, Q => Q(12)
                           , QN => n151);
   Q_reg_11_inst : DFFR_X1 port map( D => n120, CK => CK, RN => n97, Q => Q(11)
                           , QN => n152);
   Q_reg_10_inst : DFFR_X1 port map( D => n121, CK => CK, RN => n97, Q => Q(10)
                           , QN => n153);
   Q_reg_9_inst : DFFR_X1 port map( D => n122, CK => CK, RN => n97, Q => Q(9), 
                           QN => n154);
   Q_reg_8_inst : DFFR_X1 port map( D => n123, CK => CK, RN => n97, Q => Q(8), 
                           QN => n155);
   Q_reg_7_inst : DFFR_X1 port map( D => n124, CK => CK, RN => n97, Q => Q(7), 
                           QN => n156);
   Q_reg_6_inst : DFFR_X1 port map( D => n125, CK => CK, RN => n97, Q => Q(6), 
                           QN => n157);
   Q_reg_5_inst : DFFR_X1 port map( D => n126, CK => CK, RN => n97, Q => Q(5), 
                           QN => n158);
   Q_reg_4_inst : DFFR_X1 port map( D => n127, CK => CK, RN => n97, Q => Q(4), 
                           QN => n159);
   Q_reg_3_inst : DFFR_X1 port map( D => n128, CK => CK, RN => n97, Q => Q(3), 
                           QN => n160);
   Q_reg_2_inst : DFFR_X1 port map( D => n129, CK => CK, RN => n97, Q => Q(2), 
                           QN => n161);
   Q_reg_1_inst : DFFR_X1 port map( D => n130, CK => CK, RN => n97, Q => Q(1), 
                           QN => n162);
   Q_reg_0_inst : DFFR_X1 port map( D => n131, CK => CK, RN => n97, Q => Q(0), 
                           QN => n163);
   U2 : BUF_X1 port map( A => RESET, Z => n97);
   U3 : BUF_X1 port map( A => RESET, Z => n98);
   U4 : BUF_X1 port map( A => RESET, Z => n99);
   U5 : OAI21_X1 port map( B1 => n163, B2 => ENABLE, A => n195, ZN => n131);
   U6 : NAND2_X1 port map( A1 => ENABLE, A2 => D(0), ZN => n195);
   U7 : OAI21_X1 port map( B1 => n162, B2 => ENABLE, A => n194, ZN => n130);
   U8 : NAND2_X1 port map( A1 => D(1), A2 => ENABLE, ZN => n194);
   U9 : OAI21_X1 port map( B1 => n161, B2 => ENABLE, A => n193, ZN => n129);
   U10 : NAND2_X1 port map( A1 => D(2), A2 => ENABLE, ZN => n193);
   U11 : OAI21_X1 port map( B1 => n160, B2 => ENABLE, A => n192, ZN => n128);
   U12 : NAND2_X1 port map( A1 => D(3), A2 => ENABLE, ZN => n192);
   U13 : OAI21_X1 port map( B1 => n159, B2 => ENABLE, A => n191, ZN => n127);
   U14 : NAND2_X1 port map( A1 => D(4), A2 => ENABLE, ZN => n191);
   U15 : OAI21_X1 port map( B1 => n158, B2 => ENABLE, A => n190, ZN => n126);
   U16 : NAND2_X1 port map( A1 => D(5), A2 => ENABLE, ZN => n190);
   U17 : OAI21_X1 port map( B1 => n157, B2 => ENABLE, A => n189, ZN => n125);
   U18 : NAND2_X1 port map( A1 => D(6), A2 => ENABLE, ZN => n189);
   U19 : OAI21_X1 port map( B1 => n156, B2 => ENABLE, A => n188, ZN => n124);
   U20 : NAND2_X1 port map( A1 => D(7), A2 => ENABLE, ZN => n188);
   U21 : OAI21_X1 port map( B1 => n155, B2 => ENABLE, A => n187, ZN => n123);
   U22 : NAND2_X1 port map( A1 => D(8), A2 => ENABLE, ZN => n187);
   U23 : OAI21_X1 port map( B1 => n154, B2 => ENABLE, A => n186, ZN => n122);
   U24 : NAND2_X1 port map( A1 => D(9), A2 => ENABLE, ZN => n186);
   U25 : OAI21_X1 port map( B1 => n153, B2 => ENABLE, A => n185, ZN => n121);
   U26 : NAND2_X1 port map( A1 => D(10), A2 => ENABLE, ZN => n185);
   U27 : OAI21_X1 port map( B1 => n152, B2 => ENABLE, A => n184, ZN => n120);
   U28 : NAND2_X1 port map( A1 => D(11), A2 => ENABLE, ZN => n184);
   U29 : OAI21_X1 port map( B1 => n151, B2 => ENABLE, A => n183, ZN => n119);
   U30 : NAND2_X1 port map( A1 => D(12), A2 => ENABLE, ZN => n183);
   U31 : OAI21_X1 port map( B1 => n150, B2 => ENABLE, A => n182, ZN => n118);
   U32 : NAND2_X1 port map( A1 => D(13), A2 => ENABLE, ZN => n182);
   U33 : OAI21_X1 port map( B1 => n149, B2 => ENABLE, A => n181, ZN => n117);
   U34 : NAND2_X1 port map( A1 => D(14), A2 => ENABLE, ZN => n181);
   U35 : OAI21_X1 port map( B1 => n148, B2 => ENABLE, A => n180, ZN => n116);
   U36 : NAND2_X1 port map( A1 => D(15), A2 => ENABLE, ZN => n180);
   U37 : OAI21_X1 port map( B1 => n147, B2 => ENABLE, A => n179, ZN => n115);
   U38 : NAND2_X1 port map( A1 => D(16), A2 => ENABLE, ZN => n179);
   U39 : OAI21_X1 port map( B1 => n146, B2 => ENABLE, A => n178, ZN => n114);
   U40 : NAND2_X1 port map( A1 => D(17), A2 => ENABLE, ZN => n178);
   U41 : OAI21_X1 port map( B1 => n145, B2 => ENABLE, A => n177, ZN => n113);
   U42 : NAND2_X1 port map( A1 => D(18), A2 => ENABLE, ZN => n177);
   U43 : OAI21_X1 port map( B1 => n144, B2 => ENABLE, A => n176, ZN => n112);
   U44 : NAND2_X1 port map( A1 => D(19), A2 => ENABLE, ZN => n176);
   U45 : OAI21_X1 port map( B1 => n143, B2 => ENABLE, A => n175, ZN => n111);
   U46 : NAND2_X1 port map( A1 => D(20), A2 => ENABLE, ZN => n175);
   U47 : OAI21_X1 port map( B1 => n142, B2 => ENABLE, A => n174, ZN => n110);
   U48 : NAND2_X1 port map( A1 => D(21), A2 => ENABLE, ZN => n174);
   U49 : OAI21_X1 port map( B1 => n141, B2 => ENABLE, A => n173, ZN => n109);
   U50 : NAND2_X1 port map( A1 => D(22), A2 => ENABLE, ZN => n173);
   U51 : OAI21_X1 port map( B1 => n140, B2 => ENABLE, A => n172, ZN => n108);
   U52 : NAND2_X1 port map( A1 => D(23), A2 => ENABLE, ZN => n172);
   U53 : OAI21_X1 port map( B1 => n139, B2 => ENABLE, A => n171, ZN => n107);
   U54 : NAND2_X1 port map( A1 => D(24), A2 => ENABLE, ZN => n171);
   U55 : OAI21_X1 port map( B1 => n138, B2 => ENABLE, A => n170, ZN => n106);
   U56 : NAND2_X1 port map( A1 => D(25), A2 => ENABLE, ZN => n170);
   U57 : OAI21_X1 port map( B1 => n137, B2 => ENABLE, A => n169, ZN => n105);
   U58 : NAND2_X1 port map( A1 => D(26), A2 => ENABLE, ZN => n169);
   U59 : OAI21_X1 port map( B1 => n136, B2 => ENABLE, A => n168, ZN => n104);
   U60 : NAND2_X1 port map( A1 => D(27), A2 => ENABLE, ZN => n168);
   U61 : OAI21_X1 port map( B1 => n135, B2 => ENABLE, A => n167, ZN => n103);
   U62 : NAND2_X1 port map( A1 => D(28), A2 => ENABLE, ZN => n167);
   U63 : OAI21_X1 port map( B1 => n134, B2 => ENABLE, A => n166, ZN => n102);
   U64 : NAND2_X1 port map( A1 => D(29), A2 => ENABLE, ZN => n166);
   U65 : OAI21_X1 port map( B1 => n133, B2 => ENABLE, A => n165, ZN => n101);
   U66 : NAND2_X1 port map( A1 => D(30), A2 => ENABLE, ZN => n165);
   U67 : OAI21_X1 port map( B1 => n132, B2 => ENABLE, A => n164, ZN => n100);
   U68 : NAND2_X1 port map( A1 => D(31), A2 => ENABLE, ZN => n164);

end SYN_ASYNCHBEHAV;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity regFFD_NBIT32_16 is

   port( CK, RESET, ENABLE : in std_logic;  D : in std_logic_vector (31 downto 
         0);  Q : out std_logic_vector (31 downto 0));

end regFFD_NBIT32_16;

architecture SYN_ASYNCHBEHAV of regFFD_NBIT32_16 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, 
      n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, 
      n121, n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, 
      n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, 
      n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, 
      n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, 
      n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, 
      n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, 
      n193, n194, n195 : std_logic;

begin
   
   Q_reg_31_inst : DFFR_X1 port map( D => n100, CK => CK, RN => n99, Q => Q(31)
                           , QN => n132);
   Q_reg_30_inst : DFFR_X1 port map( D => n101, CK => CK, RN => n99, Q => Q(30)
                           , QN => n133);
   Q_reg_29_inst : DFFR_X1 port map( D => n102, CK => CK, RN => n99, Q => Q(29)
                           , QN => n134);
   Q_reg_28_inst : DFFR_X1 port map( D => n103, CK => CK, RN => n99, Q => Q(28)
                           , QN => n135);
   Q_reg_27_inst : DFFR_X1 port map( D => n104, CK => CK, RN => n99, Q => Q(27)
                           , QN => n136);
   Q_reg_26_inst : DFFR_X1 port map( D => n105, CK => CK, RN => n99, Q => Q(26)
                           , QN => n137);
   Q_reg_25_inst : DFFR_X1 port map( D => n106, CK => CK, RN => n99, Q => Q(25)
                           , QN => n138);
   Q_reg_24_inst : DFFR_X1 port map( D => n107, CK => CK, RN => n99, Q => Q(24)
                           , QN => n139);
   Q_reg_23_inst : DFFR_X1 port map( D => n108, CK => CK, RN => n98, Q => Q(23)
                           , QN => n140);
   Q_reg_22_inst : DFFR_X1 port map( D => n109, CK => CK, RN => n98, Q => Q(22)
                           , QN => n141);
   Q_reg_21_inst : DFFR_X1 port map( D => n110, CK => CK, RN => n98, Q => Q(21)
                           , QN => n142);
   Q_reg_20_inst : DFFR_X1 port map( D => n111, CK => CK, RN => n98, Q => Q(20)
                           , QN => n143);
   Q_reg_19_inst : DFFR_X1 port map( D => n112, CK => CK, RN => n98, Q => Q(19)
                           , QN => n144);
   Q_reg_18_inst : DFFR_X1 port map( D => n113, CK => CK, RN => n98, Q => Q(18)
                           , QN => n145);
   Q_reg_17_inst : DFFR_X1 port map( D => n114, CK => CK, RN => n98, Q => Q(17)
                           , QN => n146);
   Q_reg_16_inst : DFFR_X1 port map( D => n115, CK => CK, RN => n98, Q => Q(16)
                           , QN => n147);
   Q_reg_15_inst : DFFR_X1 port map( D => n116, CK => CK, RN => n98, Q => Q(15)
                           , QN => n148);
   Q_reg_14_inst : DFFR_X1 port map( D => n117, CK => CK, RN => n98, Q => Q(14)
                           , QN => n149);
   Q_reg_13_inst : DFFR_X1 port map( D => n118, CK => CK, RN => n98, Q => Q(13)
                           , QN => n150);
   Q_reg_12_inst : DFFR_X1 port map( D => n119, CK => CK, RN => n98, Q => Q(12)
                           , QN => n151);
   Q_reg_11_inst : DFFR_X1 port map( D => n120, CK => CK, RN => n97, Q => Q(11)
                           , QN => n152);
   Q_reg_10_inst : DFFR_X1 port map( D => n121, CK => CK, RN => n97, Q => Q(10)
                           , QN => n153);
   Q_reg_9_inst : DFFR_X1 port map( D => n122, CK => CK, RN => n97, Q => Q(9), 
                           QN => n154);
   Q_reg_8_inst : DFFR_X1 port map( D => n123, CK => CK, RN => n97, Q => Q(8), 
                           QN => n155);
   Q_reg_7_inst : DFFR_X1 port map( D => n124, CK => CK, RN => n97, Q => Q(7), 
                           QN => n156);
   Q_reg_6_inst : DFFR_X1 port map( D => n125, CK => CK, RN => n97, Q => Q(6), 
                           QN => n157);
   Q_reg_5_inst : DFFR_X1 port map( D => n126, CK => CK, RN => n97, Q => Q(5), 
                           QN => n158);
   Q_reg_4_inst : DFFR_X1 port map( D => n127, CK => CK, RN => n97, Q => Q(4), 
                           QN => n159);
   Q_reg_3_inst : DFFR_X1 port map( D => n128, CK => CK, RN => n97, Q => Q(3), 
                           QN => n160);
   Q_reg_2_inst : DFFR_X1 port map( D => n129, CK => CK, RN => n97, Q => Q(2), 
                           QN => n161);
   Q_reg_1_inst : DFFR_X1 port map( D => n130, CK => CK, RN => n97, Q => Q(1), 
                           QN => n162);
   Q_reg_0_inst : DFFR_X1 port map( D => n131, CK => CK, RN => n97, Q => Q(0), 
                           QN => n163);
   U2 : BUF_X1 port map( A => RESET, Z => n97);
   U3 : BUF_X1 port map( A => RESET, Z => n98);
   U4 : BUF_X1 port map( A => RESET, Z => n99);
   U5 : OAI21_X1 port map( B1 => n163, B2 => ENABLE, A => n195, ZN => n131);
   U6 : NAND2_X1 port map( A1 => ENABLE, A2 => D(0), ZN => n195);
   U7 : OAI21_X1 port map( B1 => n162, B2 => ENABLE, A => n194, ZN => n130);
   U8 : NAND2_X1 port map( A1 => D(1), A2 => ENABLE, ZN => n194);
   U9 : OAI21_X1 port map( B1 => n161, B2 => ENABLE, A => n193, ZN => n129);
   U10 : NAND2_X1 port map( A1 => D(2), A2 => ENABLE, ZN => n193);
   U11 : OAI21_X1 port map( B1 => n160, B2 => ENABLE, A => n192, ZN => n128);
   U12 : NAND2_X1 port map( A1 => D(3), A2 => ENABLE, ZN => n192);
   U13 : OAI21_X1 port map( B1 => n159, B2 => ENABLE, A => n191, ZN => n127);
   U14 : NAND2_X1 port map( A1 => D(4), A2 => ENABLE, ZN => n191);
   U15 : OAI21_X1 port map( B1 => n158, B2 => ENABLE, A => n190, ZN => n126);
   U16 : NAND2_X1 port map( A1 => D(5), A2 => ENABLE, ZN => n190);
   U17 : OAI21_X1 port map( B1 => n157, B2 => ENABLE, A => n189, ZN => n125);
   U18 : NAND2_X1 port map( A1 => D(6), A2 => ENABLE, ZN => n189);
   U19 : OAI21_X1 port map( B1 => n156, B2 => ENABLE, A => n188, ZN => n124);
   U20 : NAND2_X1 port map( A1 => D(7), A2 => ENABLE, ZN => n188);
   U21 : OAI21_X1 port map( B1 => n155, B2 => ENABLE, A => n187, ZN => n123);
   U22 : NAND2_X1 port map( A1 => D(8), A2 => ENABLE, ZN => n187);
   U23 : OAI21_X1 port map( B1 => n154, B2 => ENABLE, A => n186, ZN => n122);
   U24 : NAND2_X1 port map( A1 => D(9), A2 => ENABLE, ZN => n186);
   U25 : OAI21_X1 port map( B1 => n153, B2 => ENABLE, A => n185, ZN => n121);
   U26 : NAND2_X1 port map( A1 => D(10), A2 => ENABLE, ZN => n185);
   U27 : OAI21_X1 port map( B1 => n152, B2 => ENABLE, A => n184, ZN => n120);
   U28 : NAND2_X1 port map( A1 => D(11), A2 => ENABLE, ZN => n184);
   U29 : OAI21_X1 port map( B1 => n151, B2 => ENABLE, A => n183, ZN => n119);
   U30 : NAND2_X1 port map( A1 => D(12), A2 => ENABLE, ZN => n183);
   U31 : OAI21_X1 port map( B1 => n150, B2 => ENABLE, A => n182, ZN => n118);
   U32 : NAND2_X1 port map( A1 => D(13), A2 => ENABLE, ZN => n182);
   U33 : OAI21_X1 port map( B1 => n149, B2 => ENABLE, A => n181, ZN => n117);
   U34 : NAND2_X1 port map( A1 => D(14), A2 => ENABLE, ZN => n181);
   U35 : OAI21_X1 port map( B1 => n148, B2 => ENABLE, A => n180, ZN => n116);
   U36 : NAND2_X1 port map( A1 => D(15), A2 => ENABLE, ZN => n180);
   U37 : OAI21_X1 port map( B1 => n147, B2 => ENABLE, A => n179, ZN => n115);
   U38 : NAND2_X1 port map( A1 => D(16), A2 => ENABLE, ZN => n179);
   U39 : OAI21_X1 port map( B1 => n146, B2 => ENABLE, A => n178, ZN => n114);
   U40 : NAND2_X1 port map( A1 => D(17), A2 => ENABLE, ZN => n178);
   U41 : OAI21_X1 port map( B1 => n145, B2 => ENABLE, A => n177, ZN => n113);
   U42 : NAND2_X1 port map( A1 => D(18), A2 => ENABLE, ZN => n177);
   U43 : OAI21_X1 port map( B1 => n144, B2 => ENABLE, A => n176, ZN => n112);
   U44 : NAND2_X1 port map( A1 => D(19), A2 => ENABLE, ZN => n176);
   U45 : OAI21_X1 port map( B1 => n143, B2 => ENABLE, A => n175, ZN => n111);
   U46 : NAND2_X1 port map( A1 => D(20), A2 => ENABLE, ZN => n175);
   U47 : OAI21_X1 port map( B1 => n142, B2 => ENABLE, A => n174, ZN => n110);
   U48 : NAND2_X1 port map( A1 => D(21), A2 => ENABLE, ZN => n174);
   U49 : OAI21_X1 port map( B1 => n141, B2 => ENABLE, A => n173, ZN => n109);
   U50 : NAND2_X1 port map( A1 => D(22), A2 => ENABLE, ZN => n173);
   U51 : OAI21_X1 port map( B1 => n140, B2 => ENABLE, A => n172, ZN => n108);
   U52 : NAND2_X1 port map( A1 => D(23), A2 => ENABLE, ZN => n172);
   U53 : OAI21_X1 port map( B1 => n139, B2 => ENABLE, A => n171, ZN => n107);
   U54 : NAND2_X1 port map( A1 => D(24), A2 => ENABLE, ZN => n171);
   U55 : OAI21_X1 port map( B1 => n138, B2 => ENABLE, A => n170, ZN => n106);
   U56 : NAND2_X1 port map( A1 => D(25), A2 => ENABLE, ZN => n170);
   U57 : OAI21_X1 port map( B1 => n137, B2 => ENABLE, A => n169, ZN => n105);
   U58 : NAND2_X1 port map( A1 => D(26), A2 => ENABLE, ZN => n169);
   U59 : OAI21_X1 port map( B1 => n136, B2 => ENABLE, A => n168, ZN => n104);
   U60 : NAND2_X1 port map( A1 => D(27), A2 => ENABLE, ZN => n168);
   U61 : OAI21_X1 port map( B1 => n135, B2 => ENABLE, A => n167, ZN => n103);
   U62 : NAND2_X1 port map( A1 => D(28), A2 => ENABLE, ZN => n167);
   U63 : OAI21_X1 port map( B1 => n134, B2 => ENABLE, A => n166, ZN => n102);
   U64 : NAND2_X1 port map( A1 => D(29), A2 => ENABLE, ZN => n166);
   U65 : OAI21_X1 port map( B1 => n133, B2 => ENABLE, A => n165, ZN => n101);
   U66 : NAND2_X1 port map( A1 => D(30), A2 => ENABLE, ZN => n165);
   U67 : OAI21_X1 port map( B1 => n132, B2 => ENABLE, A => n164, ZN => n100);
   U68 : NAND2_X1 port map( A1 => D(31), A2 => ENABLE, ZN => n164);

end SYN_ASYNCHBEHAV;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity regFFD_NBIT32_15 is

   port( CK, RESET, ENABLE : in std_logic;  D : in std_logic_vector (31 downto 
         0);  Q : out std_logic_vector (31 downto 0));

end regFFD_NBIT32_15;

architecture SYN_ASYNCHBEHAV of regFFD_NBIT32_15 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, 
      n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, 
      n121, n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, 
      n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, 
      n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, 
      n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, 
      n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, 
      n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, 
      n193, n194, n195 : std_logic;

begin
   
   Q_reg_31_inst : DFFR_X1 port map( D => n100, CK => CK, RN => n99, Q => Q(31)
                           , QN => n132);
   Q_reg_30_inst : DFFR_X1 port map( D => n101, CK => CK, RN => n99, Q => Q(30)
                           , QN => n133);
   Q_reg_29_inst : DFFR_X1 port map( D => n102, CK => CK, RN => n99, Q => Q(29)
                           , QN => n134);
   Q_reg_28_inst : DFFR_X1 port map( D => n103, CK => CK, RN => n99, Q => Q(28)
                           , QN => n135);
   Q_reg_27_inst : DFFR_X1 port map( D => n104, CK => CK, RN => n99, Q => Q(27)
                           , QN => n136);
   Q_reg_26_inst : DFFR_X1 port map( D => n105, CK => CK, RN => n99, Q => Q(26)
                           , QN => n137);
   Q_reg_25_inst : DFFR_X1 port map( D => n106, CK => CK, RN => n99, Q => Q(25)
                           , QN => n138);
   Q_reg_24_inst : DFFR_X1 port map( D => n107, CK => CK, RN => n99, Q => Q(24)
                           , QN => n139);
   Q_reg_23_inst : DFFR_X1 port map( D => n108, CK => CK, RN => n98, Q => Q(23)
                           , QN => n140);
   Q_reg_22_inst : DFFR_X1 port map( D => n109, CK => CK, RN => n98, Q => Q(22)
                           , QN => n141);
   Q_reg_21_inst : DFFR_X1 port map( D => n110, CK => CK, RN => n98, Q => Q(21)
                           , QN => n142);
   Q_reg_20_inst : DFFR_X1 port map( D => n111, CK => CK, RN => n98, Q => Q(20)
                           , QN => n143);
   Q_reg_19_inst : DFFR_X1 port map( D => n112, CK => CK, RN => n98, Q => Q(19)
                           , QN => n144);
   Q_reg_18_inst : DFFR_X1 port map( D => n113, CK => CK, RN => n98, Q => Q(18)
                           , QN => n145);
   Q_reg_17_inst : DFFR_X1 port map( D => n114, CK => CK, RN => n98, Q => Q(17)
                           , QN => n146);
   Q_reg_16_inst : DFFR_X1 port map( D => n115, CK => CK, RN => n98, Q => Q(16)
                           , QN => n147);
   Q_reg_15_inst : DFFR_X1 port map( D => n116, CK => CK, RN => n98, Q => Q(15)
                           , QN => n148);
   Q_reg_14_inst : DFFR_X1 port map( D => n117, CK => CK, RN => n98, Q => Q(14)
                           , QN => n149);
   Q_reg_13_inst : DFFR_X1 port map( D => n118, CK => CK, RN => n98, Q => Q(13)
                           , QN => n150);
   Q_reg_12_inst : DFFR_X1 port map( D => n119, CK => CK, RN => n98, Q => Q(12)
                           , QN => n151);
   Q_reg_11_inst : DFFR_X1 port map( D => n120, CK => CK, RN => n97, Q => Q(11)
                           , QN => n152);
   Q_reg_10_inst : DFFR_X1 port map( D => n121, CK => CK, RN => n97, Q => Q(10)
                           , QN => n153);
   Q_reg_9_inst : DFFR_X1 port map( D => n122, CK => CK, RN => n97, Q => Q(9), 
                           QN => n154);
   Q_reg_8_inst : DFFR_X1 port map( D => n123, CK => CK, RN => n97, Q => Q(8), 
                           QN => n155);
   Q_reg_7_inst : DFFR_X1 port map( D => n124, CK => CK, RN => n97, Q => Q(7), 
                           QN => n156);
   Q_reg_6_inst : DFFR_X1 port map( D => n125, CK => CK, RN => n97, Q => Q(6), 
                           QN => n157);
   Q_reg_5_inst : DFFR_X1 port map( D => n126, CK => CK, RN => n97, Q => Q(5), 
                           QN => n158);
   Q_reg_4_inst : DFFR_X1 port map( D => n127, CK => CK, RN => n97, Q => Q(4), 
                           QN => n159);
   Q_reg_3_inst : DFFR_X1 port map( D => n128, CK => CK, RN => n97, Q => Q(3), 
                           QN => n160);
   Q_reg_2_inst : DFFR_X1 port map( D => n129, CK => CK, RN => n97, Q => Q(2), 
                           QN => n161);
   Q_reg_1_inst : DFFR_X1 port map( D => n130, CK => CK, RN => n97, Q => Q(1), 
                           QN => n162);
   Q_reg_0_inst : DFFR_X1 port map( D => n131, CK => CK, RN => n97, Q => Q(0), 
                           QN => n163);
   U2 : BUF_X1 port map( A => RESET, Z => n97);
   U3 : BUF_X1 port map( A => RESET, Z => n98);
   U4 : BUF_X1 port map( A => RESET, Z => n99);
   U5 : OAI21_X1 port map( B1 => n163, B2 => ENABLE, A => n195, ZN => n131);
   U6 : NAND2_X1 port map( A1 => ENABLE, A2 => D(0), ZN => n195);
   U7 : OAI21_X1 port map( B1 => n162, B2 => ENABLE, A => n194, ZN => n130);
   U8 : NAND2_X1 port map( A1 => D(1), A2 => ENABLE, ZN => n194);
   U9 : OAI21_X1 port map( B1 => n161, B2 => ENABLE, A => n193, ZN => n129);
   U10 : NAND2_X1 port map( A1 => D(2), A2 => ENABLE, ZN => n193);
   U11 : OAI21_X1 port map( B1 => n160, B2 => ENABLE, A => n192, ZN => n128);
   U12 : NAND2_X1 port map( A1 => D(3), A2 => ENABLE, ZN => n192);
   U13 : OAI21_X1 port map( B1 => n159, B2 => ENABLE, A => n191, ZN => n127);
   U14 : NAND2_X1 port map( A1 => D(4), A2 => ENABLE, ZN => n191);
   U15 : OAI21_X1 port map( B1 => n158, B2 => ENABLE, A => n190, ZN => n126);
   U16 : NAND2_X1 port map( A1 => D(5), A2 => ENABLE, ZN => n190);
   U17 : OAI21_X1 port map( B1 => n157, B2 => ENABLE, A => n189, ZN => n125);
   U18 : NAND2_X1 port map( A1 => D(6), A2 => ENABLE, ZN => n189);
   U19 : OAI21_X1 port map( B1 => n156, B2 => ENABLE, A => n188, ZN => n124);
   U20 : NAND2_X1 port map( A1 => D(7), A2 => ENABLE, ZN => n188);
   U21 : OAI21_X1 port map( B1 => n155, B2 => ENABLE, A => n187, ZN => n123);
   U22 : NAND2_X1 port map( A1 => D(8), A2 => ENABLE, ZN => n187);
   U23 : OAI21_X1 port map( B1 => n154, B2 => ENABLE, A => n186, ZN => n122);
   U24 : NAND2_X1 port map( A1 => D(9), A2 => ENABLE, ZN => n186);
   U25 : OAI21_X1 port map( B1 => n153, B2 => ENABLE, A => n185, ZN => n121);
   U26 : NAND2_X1 port map( A1 => D(10), A2 => ENABLE, ZN => n185);
   U27 : OAI21_X1 port map( B1 => n152, B2 => ENABLE, A => n184, ZN => n120);
   U28 : NAND2_X1 port map( A1 => D(11), A2 => ENABLE, ZN => n184);
   U29 : OAI21_X1 port map( B1 => n151, B2 => ENABLE, A => n183, ZN => n119);
   U30 : NAND2_X1 port map( A1 => D(12), A2 => ENABLE, ZN => n183);
   U31 : OAI21_X1 port map( B1 => n150, B2 => ENABLE, A => n182, ZN => n118);
   U32 : NAND2_X1 port map( A1 => D(13), A2 => ENABLE, ZN => n182);
   U33 : OAI21_X1 port map( B1 => n149, B2 => ENABLE, A => n181, ZN => n117);
   U34 : NAND2_X1 port map( A1 => D(14), A2 => ENABLE, ZN => n181);
   U35 : OAI21_X1 port map( B1 => n148, B2 => ENABLE, A => n180, ZN => n116);
   U36 : NAND2_X1 port map( A1 => D(15), A2 => ENABLE, ZN => n180);
   U37 : OAI21_X1 port map( B1 => n147, B2 => ENABLE, A => n179, ZN => n115);
   U38 : NAND2_X1 port map( A1 => D(16), A2 => ENABLE, ZN => n179);
   U39 : OAI21_X1 port map( B1 => n146, B2 => ENABLE, A => n178, ZN => n114);
   U40 : NAND2_X1 port map( A1 => D(17), A2 => ENABLE, ZN => n178);
   U41 : OAI21_X1 port map( B1 => n145, B2 => ENABLE, A => n177, ZN => n113);
   U42 : NAND2_X1 port map( A1 => D(18), A2 => ENABLE, ZN => n177);
   U43 : OAI21_X1 port map( B1 => n144, B2 => ENABLE, A => n176, ZN => n112);
   U44 : NAND2_X1 port map( A1 => D(19), A2 => ENABLE, ZN => n176);
   U45 : OAI21_X1 port map( B1 => n143, B2 => ENABLE, A => n175, ZN => n111);
   U46 : NAND2_X1 port map( A1 => D(20), A2 => ENABLE, ZN => n175);
   U47 : OAI21_X1 port map( B1 => n142, B2 => ENABLE, A => n174, ZN => n110);
   U48 : NAND2_X1 port map( A1 => D(21), A2 => ENABLE, ZN => n174);
   U49 : OAI21_X1 port map( B1 => n141, B2 => ENABLE, A => n173, ZN => n109);
   U50 : NAND2_X1 port map( A1 => D(22), A2 => ENABLE, ZN => n173);
   U51 : OAI21_X1 port map( B1 => n140, B2 => ENABLE, A => n172, ZN => n108);
   U52 : NAND2_X1 port map( A1 => D(23), A2 => ENABLE, ZN => n172);
   U53 : OAI21_X1 port map( B1 => n139, B2 => ENABLE, A => n171, ZN => n107);
   U54 : NAND2_X1 port map( A1 => D(24), A2 => ENABLE, ZN => n171);
   U55 : OAI21_X1 port map( B1 => n138, B2 => ENABLE, A => n170, ZN => n106);
   U56 : NAND2_X1 port map( A1 => D(25), A2 => ENABLE, ZN => n170);
   U57 : OAI21_X1 port map( B1 => n137, B2 => ENABLE, A => n169, ZN => n105);
   U58 : NAND2_X1 port map( A1 => D(26), A2 => ENABLE, ZN => n169);
   U59 : OAI21_X1 port map( B1 => n136, B2 => ENABLE, A => n168, ZN => n104);
   U60 : NAND2_X1 port map( A1 => D(27), A2 => ENABLE, ZN => n168);
   U61 : OAI21_X1 port map( B1 => n135, B2 => ENABLE, A => n167, ZN => n103);
   U62 : NAND2_X1 port map( A1 => D(28), A2 => ENABLE, ZN => n167);
   U63 : OAI21_X1 port map( B1 => n134, B2 => ENABLE, A => n166, ZN => n102);
   U64 : NAND2_X1 port map( A1 => D(29), A2 => ENABLE, ZN => n166);
   U65 : OAI21_X1 port map( B1 => n133, B2 => ENABLE, A => n165, ZN => n101);
   U66 : NAND2_X1 port map( A1 => D(30), A2 => ENABLE, ZN => n165);
   U67 : OAI21_X1 port map( B1 => n132, B2 => ENABLE, A => n164, ZN => n100);
   U68 : NAND2_X1 port map( A1 => D(31), A2 => ENABLE, ZN => n164);

end SYN_ASYNCHBEHAV;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity regFFD_NBIT32_14 is

   port( CK, RESET, ENABLE : in std_logic;  D : in std_logic_vector (31 downto 
         0);  Q : out std_logic_vector (31 downto 0));

end regFFD_NBIT32_14;

architecture SYN_ASYNCHBEHAV of regFFD_NBIT32_14 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, 
      n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, 
      n121, n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, 
      n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, 
      n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, 
      n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, 
      n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, 
      n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, 
      n193, n194, n195 : std_logic;

begin
   
   Q_reg_31_inst : DFFR_X1 port map( D => n100, CK => CK, RN => n99, Q => Q(31)
                           , QN => n132);
   Q_reg_30_inst : DFFR_X1 port map( D => n101, CK => CK, RN => n99, Q => Q(30)
                           , QN => n133);
   Q_reg_29_inst : DFFR_X1 port map( D => n102, CK => CK, RN => n99, Q => Q(29)
                           , QN => n134);
   Q_reg_28_inst : DFFR_X1 port map( D => n103, CK => CK, RN => n99, Q => Q(28)
                           , QN => n135);
   Q_reg_27_inst : DFFR_X1 port map( D => n104, CK => CK, RN => n99, Q => Q(27)
                           , QN => n136);
   Q_reg_26_inst : DFFR_X1 port map( D => n105, CK => CK, RN => n99, Q => Q(26)
                           , QN => n137);
   Q_reg_25_inst : DFFR_X1 port map( D => n106, CK => CK, RN => n99, Q => Q(25)
                           , QN => n138);
   Q_reg_24_inst : DFFR_X1 port map( D => n107, CK => CK, RN => n99, Q => Q(24)
                           , QN => n139);
   Q_reg_23_inst : DFFR_X1 port map( D => n108, CK => CK, RN => n98, Q => Q(23)
                           , QN => n140);
   Q_reg_22_inst : DFFR_X1 port map( D => n109, CK => CK, RN => n98, Q => Q(22)
                           , QN => n141);
   Q_reg_21_inst : DFFR_X1 port map( D => n110, CK => CK, RN => n98, Q => Q(21)
                           , QN => n142);
   Q_reg_20_inst : DFFR_X1 port map( D => n111, CK => CK, RN => n98, Q => Q(20)
                           , QN => n143);
   Q_reg_19_inst : DFFR_X1 port map( D => n112, CK => CK, RN => n98, Q => Q(19)
                           , QN => n144);
   Q_reg_18_inst : DFFR_X1 port map( D => n113, CK => CK, RN => n98, Q => Q(18)
                           , QN => n145);
   Q_reg_17_inst : DFFR_X1 port map( D => n114, CK => CK, RN => n98, Q => Q(17)
                           , QN => n146);
   Q_reg_16_inst : DFFR_X1 port map( D => n115, CK => CK, RN => n98, Q => Q(16)
                           , QN => n147);
   Q_reg_15_inst : DFFR_X1 port map( D => n116, CK => CK, RN => n98, Q => Q(15)
                           , QN => n148);
   Q_reg_14_inst : DFFR_X1 port map( D => n117, CK => CK, RN => n98, Q => Q(14)
                           , QN => n149);
   Q_reg_13_inst : DFFR_X1 port map( D => n118, CK => CK, RN => n98, Q => Q(13)
                           , QN => n150);
   Q_reg_12_inst : DFFR_X1 port map( D => n119, CK => CK, RN => n98, Q => Q(12)
                           , QN => n151);
   Q_reg_11_inst : DFFR_X1 port map( D => n120, CK => CK, RN => n97, Q => Q(11)
                           , QN => n152);
   Q_reg_10_inst : DFFR_X1 port map( D => n121, CK => CK, RN => n97, Q => Q(10)
                           , QN => n153);
   Q_reg_9_inst : DFFR_X1 port map( D => n122, CK => CK, RN => n97, Q => Q(9), 
                           QN => n154);
   Q_reg_8_inst : DFFR_X1 port map( D => n123, CK => CK, RN => n97, Q => Q(8), 
                           QN => n155);
   Q_reg_7_inst : DFFR_X1 port map( D => n124, CK => CK, RN => n97, Q => Q(7), 
                           QN => n156);
   Q_reg_6_inst : DFFR_X1 port map( D => n125, CK => CK, RN => n97, Q => Q(6), 
                           QN => n157);
   Q_reg_5_inst : DFFR_X1 port map( D => n126, CK => CK, RN => n97, Q => Q(5), 
                           QN => n158);
   Q_reg_4_inst : DFFR_X1 port map( D => n127, CK => CK, RN => n97, Q => Q(4), 
                           QN => n159);
   Q_reg_3_inst : DFFR_X1 port map( D => n128, CK => CK, RN => n97, Q => Q(3), 
                           QN => n160);
   Q_reg_2_inst : DFFR_X1 port map( D => n129, CK => CK, RN => n97, Q => Q(2), 
                           QN => n161);
   Q_reg_1_inst : DFFR_X1 port map( D => n130, CK => CK, RN => n97, Q => Q(1), 
                           QN => n162);
   Q_reg_0_inst : DFFR_X1 port map( D => n131, CK => CK, RN => n97, Q => Q(0), 
                           QN => n163);
   U2 : BUF_X1 port map( A => RESET, Z => n97);
   U3 : BUF_X1 port map( A => RESET, Z => n98);
   U4 : BUF_X1 port map( A => RESET, Z => n99);
   U5 : OAI21_X1 port map( B1 => n163, B2 => ENABLE, A => n195, ZN => n131);
   U6 : NAND2_X1 port map( A1 => ENABLE, A2 => D(0), ZN => n195);
   U7 : OAI21_X1 port map( B1 => n162, B2 => ENABLE, A => n194, ZN => n130);
   U8 : NAND2_X1 port map( A1 => D(1), A2 => ENABLE, ZN => n194);
   U9 : OAI21_X1 port map( B1 => n161, B2 => ENABLE, A => n193, ZN => n129);
   U10 : NAND2_X1 port map( A1 => D(2), A2 => ENABLE, ZN => n193);
   U11 : OAI21_X1 port map( B1 => n160, B2 => ENABLE, A => n192, ZN => n128);
   U12 : NAND2_X1 port map( A1 => D(3), A2 => ENABLE, ZN => n192);
   U13 : OAI21_X1 port map( B1 => n159, B2 => ENABLE, A => n191, ZN => n127);
   U14 : NAND2_X1 port map( A1 => D(4), A2 => ENABLE, ZN => n191);
   U15 : OAI21_X1 port map( B1 => n158, B2 => ENABLE, A => n190, ZN => n126);
   U16 : NAND2_X1 port map( A1 => D(5), A2 => ENABLE, ZN => n190);
   U17 : OAI21_X1 port map( B1 => n157, B2 => ENABLE, A => n189, ZN => n125);
   U18 : NAND2_X1 port map( A1 => D(6), A2 => ENABLE, ZN => n189);
   U19 : OAI21_X1 port map( B1 => n156, B2 => ENABLE, A => n188, ZN => n124);
   U20 : NAND2_X1 port map( A1 => D(7), A2 => ENABLE, ZN => n188);
   U21 : OAI21_X1 port map( B1 => n155, B2 => ENABLE, A => n187, ZN => n123);
   U22 : NAND2_X1 port map( A1 => D(8), A2 => ENABLE, ZN => n187);
   U23 : OAI21_X1 port map( B1 => n154, B2 => ENABLE, A => n186, ZN => n122);
   U24 : NAND2_X1 port map( A1 => D(9), A2 => ENABLE, ZN => n186);
   U25 : OAI21_X1 port map( B1 => n153, B2 => ENABLE, A => n185, ZN => n121);
   U26 : NAND2_X1 port map( A1 => D(10), A2 => ENABLE, ZN => n185);
   U27 : OAI21_X1 port map( B1 => n152, B2 => ENABLE, A => n184, ZN => n120);
   U28 : NAND2_X1 port map( A1 => D(11), A2 => ENABLE, ZN => n184);
   U29 : OAI21_X1 port map( B1 => n151, B2 => ENABLE, A => n183, ZN => n119);
   U30 : NAND2_X1 port map( A1 => D(12), A2 => ENABLE, ZN => n183);
   U31 : OAI21_X1 port map( B1 => n150, B2 => ENABLE, A => n182, ZN => n118);
   U32 : NAND2_X1 port map( A1 => D(13), A2 => ENABLE, ZN => n182);
   U33 : OAI21_X1 port map( B1 => n149, B2 => ENABLE, A => n181, ZN => n117);
   U34 : NAND2_X1 port map( A1 => D(14), A2 => ENABLE, ZN => n181);
   U35 : OAI21_X1 port map( B1 => n148, B2 => ENABLE, A => n180, ZN => n116);
   U36 : NAND2_X1 port map( A1 => D(15), A2 => ENABLE, ZN => n180);
   U37 : OAI21_X1 port map( B1 => n147, B2 => ENABLE, A => n179, ZN => n115);
   U38 : NAND2_X1 port map( A1 => D(16), A2 => ENABLE, ZN => n179);
   U39 : OAI21_X1 port map( B1 => n146, B2 => ENABLE, A => n178, ZN => n114);
   U40 : NAND2_X1 port map( A1 => D(17), A2 => ENABLE, ZN => n178);
   U41 : OAI21_X1 port map( B1 => n145, B2 => ENABLE, A => n177, ZN => n113);
   U42 : NAND2_X1 port map( A1 => D(18), A2 => ENABLE, ZN => n177);
   U43 : OAI21_X1 port map( B1 => n144, B2 => ENABLE, A => n176, ZN => n112);
   U44 : NAND2_X1 port map( A1 => D(19), A2 => ENABLE, ZN => n176);
   U45 : OAI21_X1 port map( B1 => n143, B2 => ENABLE, A => n175, ZN => n111);
   U46 : NAND2_X1 port map( A1 => D(20), A2 => ENABLE, ZN => n175);
   U47 : OAI21_X1 port map( B1 => n142, B2 => ENABLE, A => n174, ZN => n110);
   U48 : NAND2_X1 port map( A1 => D(21), A2 => ENABLE, ZN => n174);
   U49 : OAI21_X1 port map( B1 => n141, B2 => ENABLE, A => n173, ZN => n109);
   U50 : NAND2_X1 port map( A1 => D(22), A2 => ENABLE, ZN => n173);
   U51 : OAI21_X1 port map( B1 => n140, B2 => ENABLE, A => n172, ZN => n108);
   U52 : NAND2_X1 port map( A1 => D(23), A2 => ENABLE, ZN => n172);
   U53 : OAI21_X1 port map( B1 => n139, B2 => ENABLE, A => n171, ZN => n107);
   U54 : NAND2_X1 port map( A1 => D(24), A2 => ENABLE, ZN => n171);
   U55 : OAI21_X1 port map( B1 => n138, B2 => ENABLE, A => n170, ZN => n106);
   U56 : NAND2_X1 port map( A1 => D(25), A2 => ENABLE, ZN => n170);
   U57 : OAI21_X1 port map( B1 => n137, B2 => ENABLE, A => n169, ZN => n105);
   U58 : NAND2_X1 port map( A1 => D(26), A2 => ENABLE, ZN => n169);
   U59 : OAI21_X1 port map( B1 => n136, B2 => ENABLE, A => n168, ZN => n104);
   U60 : NAND2_X1 port map( A1 => D(27), A2 => ENABLE, ZN => n168);
   U61 : OAI21_X1 port map( B1 => n135, B2 => ENABLE, A => n167, ZN => n103);
   U62 : NAND2_X1 port map( A1 => D(28), A2 => ENABLE, ZN => n167);
   U63 : OAI21_X1 port map( B1 => n134, B2 => ENABLE, A => n166, ZN => n102);
   U64 : NAND2_X1 port map( A1 => D(29), A2 => ENABLE, ZN => n166);
   U65 : OAI21_X1 port map( B1 => n133, B2 => ENABLE, A => n165, ZN => n101);
   U66 : NAND2_X1 port map( A1 => D(30), A2 => ENABLE, ZN => n165);
   U67 : OAI21_X1 port map( B1 => n132, B2 => ENABLE, A => n164, ZN => n100);
   U68 : NAND2_X1 port map( A1 => D(31), A2 => ENABLE, ZN => n164);

end SYN_ASYNCHBEHAV;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity regFFD_NBIT32_13 is

   port( CK, RESET, ENABLE : in std_logic;  D : in std_logic_vector (31 downto 
         0);  Q : out std_logic_vector (31 downto 0));

end regFFD_NBIT32_13;

architecture SYN_ASYNCHBEHAV of regFFD_NBIT32_13 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, 
      n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, 
      n121, n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, 
      n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, 
      n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, 
      n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, 
      n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, 
      n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, 
      n193, n194, n195 : std_logic;

begin
   
   Q_reg_31_inst : DFFR_X1 port map( D => n100, CK => CK, RN => n99, Q => Q(31)
                           , QN => n132);
   Q_reg_30_inst : DFFR_X1 port map( D => n101, CK => CK, RN => n99, Q => Q(30)
                           , QN => n133);
   Q_reg_29_inst : DFFR_X1 port map( D => n102, CK => CK, RN => n99, Q => Q(29)
                           , QN => n134);
   Q_reg_28_inst : DFFR_X1 port map( D => n103, CK => CK, RN => n99, Q => Q(28)
                           , QN => n135);
   Q_reg_27_inst : DFFR_X1 port map( D => n104, CK => CK, RN => n99, Q => Q(27)
                           , QN => n136);
   Q_reg_26_inst : DFFR_X1 port map( D => n105, CK => CK, RN => n99, Q => Q(26)
                           , QN => n137);
   Q_reg_25_inst : DFFR_X1 port map( D => n106, CK => CK, RN => n99, Q => Q(25)
                           , QN => n138);
   Q_reg_24_inst : DFFR_X1 port map( D => n107, CK => CK, RN => n99, Q => Q(24)
                           , QN => n139);
   Q_reg_23_inst : DFFR_X1 port map( D => n108, CK => CK, RN => n98, Q => Q(23)
                           , QN => n140);
   Q_reg_22_inst : DFFR_X1 port map( D => n109, CK => CK, RN => n98, Q => Q(22)
                           , QN => n141);
   Q_reg_21_inst : DFFR_X1 port map( D => n110, CK => CK, RN => n98, Q => Q(21)
                           , QN => n142);
   Q_reg_20_inst : DFFR_X1 port map( D => n111, CK => CK, RN => n98, Q => Q(20)
                           , QN => n143);
   Q_reg_19_inst : DFFR_X1 port map( D => n112, CK => CK, RN => n98, Q => Q(19)
                           , QN => n144);
   Q_reg_18_inst : DFFR_X1 port map( D => n113, CK => CK, RN => n98, Q => Q(18)
                           , QN => n145);
   Q_reg_17_inst : DFFR_X1 port map( D => n114, CK => CK, RN => n98, Q => Q(17)
                           , QN => n146);
   Q_reg_16_inst : DFFR_X1 port map( D => n115, CK => CK, RN => n98, Q => Q(16)
                           , QN => n147);
   Q_reg_15_inst : DFFR_X1 port map( D => n116, CK => CK, RN => n98, Q => Q(15)
                           , QN => n148);
   Q_reg_14_inst : DFFR_X1 port map( D => n117, CK => CK, RN => n98, Q => Q(14)
                           , QN => n149);
   Q_reg_13_inst : DFFR_X1 port map( D => n118, CK => CK, RN => n98, Q => Q(13)
                           , QN => n150);
   Q_reg_12_inst : DFFR_X1 port map( D => n119, CK => CK, RN => n98, Q => Q(12)
                           , QN => n151);
   Q_reg_11_inst : DFFR_X1 port map( D => n120, CK => CK, RN => n97, Q => Q(11)
                           , QN => n152);
   Q_reg_10_inst : DFFR_X1 port map( D => n121, CK => CK, RN => n97, Q => Q(10)
                           , QN => n153);
   Q_reg_9_inst : DFFR_X1 port map( D => n122, CK => CK, RN => n97, Q => Q(9), 
                           QN => n154);
   Q_reg_8_inst : DFFR_X1 port map( D => n123, CK => CK, RN => n97, Q => Q(8), 
                           QN => n155);
   Q_reg_7_inst : DFFR_X1 port map( D => n124, CK => CK, RN => n97, Q => Q(7), 
                           QN => n156);
   Q_reg_6_inst : DFFR_X1 port map( D => n125, CK => CK, RN => n97, Q => Q(6), 
                           QN => n157);
   Q_reg_5_inst : DFFR_X1 port map( D => n126, CK => CK, RN => n97, Q => Q(5), 
                           QN => n158);
   Q_reg_4_inst : DFFR_X1 port map( D => n127, CK => CK, RN => n97, Q => Q(4), 
                           QN => n159);
   Q_reg_3_inst : DFFR_X1 port map( D => n128, CK => CK, RN => n97, Q => Q(3), 
                           QN => n160);
   Q_reg_2_inst : DFFR_X1 port map( D => n129, CK => CK, RN => n97, Q => Q(2), 
                           QN => n161);
   Q_reg_1_inst : DFFR_X1 port map( D => n130, CK => CK, RN => n97, Q => Q(1), 
                           QN => n162);
   Q_reg_0_inst : DFFR_X1 port map( D => n131, CK => CK, RN => n97, Q => Q(0), 
                           QN => n163);
   U2 : BUF_X1 port map( A => RESET, Z => n97);
   U3 : BUF_X1 port map( A => RESET, Z => n98);
   U4 : BUF_X1 port map( A => RESET, Z => n99);
   U5 : OAI21_X1 port map( B1 => n163, B2 => ENABLE, A => n195, ZN => n131);
   U6 : NAND2_X1 port map( A1 => ENABLE, A2 => D(0), ZN => n195);
   U7 : OAI21_X1 port map( B1 => n162, B2 => ENABLE, A => n194, ZN => n130);
   U8 : NAND2_X1 port map( A1 => D(1), A2 => ENABLE, ZN => n194);
   U9 : OAI21_X1 port map( B1 => n161, B2 => ENABLE, A => n193, ZN => n129);
   U10 : NAND2_X1 port map( A1 => D(2), A2 => ENABLE, ZN => n193);
   U11 : OAI21_X1 port map( B1 => n160, B2 => ENABLE, A => n192, ZN => n128);
   U12 : NAND2_X1 port map( A1 => D(3), A2 => ENABLE, ZN => n192);
   U13 : OAI21_X1 port map( B1 => n159, B2 => ENABLE, A => n191, ZN => n127);
   U14 : NAND2_X1 port map( A1 => D(4), A2 => ENABLE, ZN => n191);
   U15 : OAI21_X1 port map( B1 => n158, B2 => ENABLE, A => n190, ZN => n126);
   U16 : NAND2_X1 port map( A1 => D(5), A2 => ENABLE, ZN => n190);
   U17 : OAI21_X1 port map( B1 => n157, B2 => ENABLE, A => n189, ZN => n125);
   U18 : NAND2_X1 port map( A1 => D(6), A2 => ENABLE, ZN => n189);
   U19 : OAI21_X1 port map( B1 => n156, B2 => ENABLE, A => n188, ZN => n124);
   U20 : NAND2_X1 port map( A1 => D(7), A2 => ENABLE, ZN => n188);
   U21 : OAI21_X1 port map( B1 => n155, B2 => ENABLE, A => n187, ZN => n123);
   U22 : NAND2_X1 port map( A1 => D(8), A2 => ENABLE, ZN => n187);
   U23 : OAI21_X1 port map( B1 => n154, B2 => ENABLE, A => n186, ZN => n122);
   U24 : NAND2_X1 port map( A1 => D(9), A2 => ENABLE, ZN => n186);
   U25 : OAI21_X1 port map( B1 => n153, B2 => ENABLE, A => n185, ZN => n121);
   U26 : NAND2_X1 port map( A1 => D(10), A2 => ENABLE, ZN => n185);
   U27 : OAI21_X1 port map( B1 => n152, B2 => ENABLE, A => n184, ZN => n120);
   U28 : NAND2_X1 port map( A1 => D(11), A2 => ENABLE, ZN => n184);
   U29 : OAI21_X1 port map( B1 => n151, B2 => ENABLE, A => n183, ZN => n119);
   U30 : NAND2_X1 port map( A1 => D(12), A2 => ENABLE, ZN => n183);
   U31 : OAI21_X1 port map( B1 => n150, B2 => ENABLE, A => n182, ZN => n118);
   U32 : NAND2_X1 port map( A1 => D(13), A2 => ENABLE, ZN => n182);
   U33 : OAI21_X1 port map( B1 => n149, B2 => ENABLE, A => n181, ZN => n117);
   U34 : NAND2_X1 port map( A1 => D(14), A2 => ENABLE, ZN => n181);
   U35 : OAI21_X1 port map( B1 => n148, B2 => ENABLE, A => n180, ZN => n116);
   U36 : NAND2_X1 port map( A1 => D(15), A2 => ENABLE, ZN => n180);
   U37 : OAI21_X1 port map( B1 => n147, B2 => ENABLE, A => n179, ZN => n115);
   U38 : NAND2_X1 port map( A1 => D(16), A2 => ENABLE, ZN => n179);
   U39 : OAI21_X1 port map( B1 => n146, B2 => ENABLE, A => n178, ZN => n114);
   U40 : NAND2_X1 port map( A1 => D(17), A2 => ENABLE, ZN => n178);
   U41 : OAI21_X1 port map( B1 => n145, B2 => ENABLE, A => n177, ZN => n113);
   U42 : NAND2_X1 port map( A1 => D(18), A2 => ENABLE, ZN => n177);
   U43 : OAI21_X1 port map( B1 => n144, B2 => ENABLE, A => n176, ZN => n112);
   U44 : NAND2_X1 port map( A1 => D(19), A2 => ENABLE, ZN => n176);
   U45 : OAI21_X1 port map( B1 => n143, B2 => ENABLE, A => n175, ZN => n111);
   U46 : NAND2_X1 port map( A1 => D(20), A2 => ENABLE, ZN => n175);
   U47 : OAI21_X1 port map( B1 => n142, B2 => ENABLE, A => n174, ZN => n110);
   U48 : NAND2_X1 port map( A1 => D(21), A2 => ENABLE, ZN => n174);
   U49 : OAI21_X1 port map( B1 => n141, B2 => ENABLE, A => n173, ZN => n109);
   U50 : NAND2_X1 port map( A1 => D(22), A2 => ENABLE, ZN => n173);
   U51 : OAI21_X1 port map( B1 => n140, B2 => ENABLE, A => n172, ZN => n108);
   U52 : NAND2_X1 port map( A1 => D(23), A2 => ENABLE, ZN => n172);
   U53 : OAI21_X1 port map( B1 => n139, B2 => ENABLE, A => n171, ZN => n107);
   U54 : NAND2_X1 port map( A1 => D(24), A2 => ENABLE, ZN => n171);
   U55 : OAI21_X1 port map( B1 => n138, B2 => ENABLE, A => n170, ZN => n106);
   U56 : NAND2_X1 port map( A1 => D(25), A2 => ENABLE, ZN => n170);
   U57 : OAI21_X1 port map( B1 => n137, B2 => ENABLE, A => n169, ZN => n105);
   U58 : NAND2_X1 port map( A1 => D(26), A2 => ENABLE, ZN => n169);
   U59 : OAI21_X1 port map( B1 => n136, B2 => ENABLE, A => n168, ZN => n104);
   U60 : NAND2_X1 port map( A1 => D(27), A2 => ENABLE, ZN => n168);
   U61 : OAI21_X1 port map( B1 => n135, B2 => ENABLE, A => n167, ZN => n103);
   U62 : NAND2_X1 port map( A1 => D(28), A2 => ENABLE, ZN => n167);
   U63 : OAI21_X1 port map( B1 => n134, B2 => ENABLE, A => n166, ZN => n102);
   U64 : NAND2_X1 port map( A1 => D(29), A2 => ENABLE, ZN => n166);
   U65 : OAI21_X1 port map( B1 => n133, B2 => ENABLE, A => n165, ZN => n101);
   U66 : NAND2_X1 port map( A1 => D(30), A2 => ENABLE, ZN => n165);
   U67 : OAI21_X1 port map( B1 => n132, B2 => ENABLE, A => n164, ZN => n100);
   U68 : NAND2_X1 port map( A1 => D(31), A2 => ENABLE, ZN => n164);

end SYN_ASYNCHBEHAV;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity regFFD_NBIT32_12 is

   port( CK, RESET, ENABLE : in std_logic;  D : in std_logic_vector (31 downto 
         0);  Q : out std_logic_vector (31 downto 0));

end regFFD_NBIT32_12;

architecture SYN_ASYNCHBEHAV of regFFD_NBIT32_12 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, 
      n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, 
      n121, n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, 
      n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, 
      n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, 
      n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, 
      n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, 
      n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, 
      n193, n194, n195 : std_logic;

begin
   
   Q_reg_31_inst : DFFR_X1 port map( D => n100, CK => CK, RN => n99, Q => Q(31)
                           , QN => n132);
   Q_reg_30_inst : DFFR_X1 port map( D => n101, CK => CK, RN => n99, Q => Q(30)
                           , QN => n133);
   Q_reg_29_inst : DFFR_X1 port map( D => n102, CK => CK, RN => n99, Q => Q(29)
                           , QN => n134);
   Q_reg_28_inst : DFFR_X1 port map( D => n103, CK => CK, RN => n99, Q => Q(28)
                           , QN => n135);
   Q_reg_27_inst : DFFR_X1 port map( D => n104, CK => CK, RN => n99, Q => Q(27)
                           , QN => n136);
   Q_reg_26_inst : DFFR_X1 port map( D => n105, CK => CK, RN => n99, Q => Q(26)
                           , QN => n137);
   Q_reg_25_inst : DFFR_X1 port map( D => n106, CK => CK, RN => n99, Q => Q(25)
                           , QN => n138);
   Q_reg_24_inst : DFFR_X1 port map( D => n107, CK => CK, RN => n99, Q => Q(24)
                           , QN => n139);
   Q_reg_23_inst : DFFR_X1 port map( D => n108, CK => CK, RN => n98, Q => Q(23)
                           , QN => n140);
   Q_reg_22_inst : DFFR_X1 port map( D => n109, CK => CK, RN => n98, Q => Q(22)
                           , QN => n141);
   Q_reg_21_inst : DFFR_X1 port map( D => n110, CK => CK, RN => n98, Q => Q(21)
                           , QN => n142);
   Q_reg_20_inst : DFFR_X1 port map( D => n111, CK => CK, RN => n98, Q => Q(20)
                           , QN => n143);
   Q_reg_19_inst : DFFR_X1 port map( D => n112, CK => CK, RN => n98, Q => Q(19)
                           , QN => n144);
   Q_reg_18_inst : DFFR_X1 port map( D => n113, CK => CK, RN => n98, Q => Q(18)
                           , QN => n145);
   Q_reg_17_inst : DFFR_X1 port map( D => n114, CK => CK, RN => n98, Q => Q(17)
                           , QN => n146);
   Q_reg_16_inst : DFFR_X1 port map( D => n115, CK => CK, RN => n98, Q => Q(16)
                           , QN => n147);
   Q_reg_15_inst : DFFR_X1 port map( D => n116, CK => CK, RN => n98, Q => Q(15)
                           , QN => n148);
   Q_reg_14_inst : DFFR_X1 port map( D => n117, CK => CK, RN => n98, Q => Q(14)
                           , QN => n149);
   Q_reg_13_inst : DFFR_X1 port map( D => n118, CK => CK, RN => n98, Q => Q(13)
                           , QN => n150);
   Q_reg_12_inst : DFFR_X1 port map( D => n119, CK => CK, RN => n98, Q => Q(12)
                           , QN => n151);
   Q_reg_11_inst : DFFR_X1 port map( D => n120, CK => CK, RN => n97, Q => Q(11)
                           , QN => n152);
   Q_reg_10_inst : DFFR_X1 port map( D => n121, CK => CK, RN => n97, Q => Q(10)
                           , QN => n153);
   Q_reg_9_inst : DFFR_X1 port map( D => n122, CK => CK, RN => n97, Q => Q(9), 
                           QN => n154);
   Q_reg_8_inst : DFFR_X1 port map( D => n123, CK => CK, RN => n97, Q => Q(8), 
                           QN => n155);
   Q_reg_7_inst : DFFR_X1 port map( D => n124, CK => CK, RN => n97, Q => Q(7), 
                           QN => n156);
   Q_reg_6_inst : DFFR_X1 port map( D => n125, CK => CK, RN => n97, Q => Q(6), 
                           QN => n157);
   Q_reg_5_inst : DFFR_X1 port map( D => n126, CK => CK, RN => n97, Q => Q(5), 
                           QN => n158);
   Q_reg_4_inst : DFFR_X1 port map( D => n127, CK => CK, RN => n97, Q => Q(4), 
                           QN => n159);
   Q_reg_3_inst : DFFR_X1 port map( D => n128, CK => CK, RN => n97, Q => Q(3), 
                           QN => n160);
   Q_reg_2_inst : DFFR_X1 port map( D => n129, CK => CK, RN => n97, Q => Q(2), 
                           QN => n161);
   Q_reg_1_inst : DFFR_X1 port map( D => n130, CK => CK, RN => n97, Q => Q(1), 
                           QN => n162);
   Q_reg_0_inst : DFFR_X1 port map( D => n131, CK => CK, RN => n97, Q => Q(0), 
                           QN => n163);
   U2 : BUF_X1 port map( A => RESET, Z => n97);
   U3 : BUF_X1 port map( A => RESET, Z => n98);
   U4 : BUF_X1 port map( A => RESET, Z => n99);
   U5 : OAI21_X1 port map( B1 => n163, B2 => ENABLE, A => n195, ZN => n131);
   U6 : NAND2_X1 port map( A1 => ENABLE, A2 => D(0), ZN => n195);
   U7 : OAI21_X1 port map( B1 => n162, B2 => ENABLE, A => n194, ZN => n130);
   U8 : NAND2_X1 port map( A1 => D(1), A2 => ENABLE, ZN => n194);
   U9 : OAI21_X1 port map( B1 => n161, B2 => ENABLE, A => n193, ZN => n129);
   U10 : NAND2_X1 port map( A1 => D(2), A2 => ENABLE, ZN => n193);
   U11 : OAI21_X1 port map( B1 => n160, B2 => ENABLE, A => n192, ZN => n128);
   U12 : NAND2_X1 port map( A1 => D(3), A2 => ENABLE, ZN => n192);
   U13 : OAI21_X1 port map( B1 => n159, B2 => ENABLE, A => n191, ZN => n127);
   U14 : NAND2_X1 port map( A1 => D(4), A2 => ENABLE, ZN => n191);
   U15 : OAI21_X1 port map( B1 => n158, B2 => ENABLE, A => n190, ZN => n126);
   U16 : NAND2_X1 port map( A1 => D(5), A2 => ENABLE, ZN => n190);
   U17 : OAI21_X1 port map( B1 => n157, B2 => ENABLE, A => n189, ZN => n125);
   U18 : NAND2_X1 port map( A1 => D(6), A2 => ENABLE, ZN => n189);
   U19 : OAI21_X1 port map( B1 => n156, B2 => ENABLE, A => n188, ZN => n124);
   U20 : NAND2_X1 port map( A1 => D(7), A2 => ENABLE, ZN => n188);
   U21 : OAI21_X1 port map( B1 => n155, B2 => ENABLE, A => n187, ZN => n123);
   U22 : NAND2_X1 port map( A1 => D(8), A2 => ENABLE, ZN => n187);
   U23 : OAI21_X1 port map( B1 => n154, B2 => ENABLE, A => n186, ZN => n122);
   U24 : NAND2_X1 port map( A1 => D(9), A2 => ENABLE, ZN => n186);
   U25 : OAI21_X1 port map( B1 => n153, B2 => ENABLE, A => n185, ZN => n121);
   U26 : NAND2_X1 port map( A1 => D(10), A2 => ENABLE, ZN => n185);
   U27 : OAI21_X1 port map( B1 => n152, B2 => ENABLE, A => n184, ZN => n120);
   U28 : NAND2_X1 port map( A1 => D(11), A2 => ENABLE, ZN => n184);
   U29 : OAI21_X1 port map( B1 => n151, B2 => ENABLE, A => n183, ZN => n119);
   U30 : NAND2_X1 port map( A1 => D(12), A2 => ENABLE, ZN => n183);
   U31 : OAI21_X1 port map( B1 => n150, B2 => ENABLE, A => n182, ZN => n118);
   U32 : NAND2_X1 port map( A1 => D(13), A2 => ENABLE, ZN => n182);
   U33 : OAI21_X1 port map( B1 => n149, B2 => ENABLE, A => n181, ZN => n117);
   U34 : NAND2_X1 port map( A1 => D(14), A2 => ENABLE, ZN => n181);
   U35 : OAI21_X1 port map( B1 => n148, B2 => ENABLE, A => n180, ZN => n116);
   U36 : NAND2_X1 port map( A1 => D(15), A2 => ENABLE, ZN => n180);
   U37 : OAI21_X1 port map( B1 => n147, B2 => ENABLE, A => n179, ZN => n115);
   U38 : NAND2_X1 port map( A1 => D(16), A2 => ENABLE, ZN => n179);
   U39 : OAI21_X1 port map( B1 => n146, B2 => ENABLE, A => n178, ZN => n114);
   U40 : NAND2_X1 port map( A1 => D(17), A2 => ENABLE, ZN => n178);
   U41 : OAI21_X1 port map( B1 => n145, B2 => ENABLE, A => n177, ZN => n113);
   U42 : NAND2_X1 port map( A1 => D(18), A2 => ENABLE, ZN => n177);
   U43 : OAI21_X1 port map( B1 => n144, B2 => ENABLE, A => n176, ZN => n112);
   U44 : NAND2_X1 port map( A1 => D(19), A2 => ENABLE, ZN => n176);
   U45 : OAI21_X1 port map( B1 => n143, B2 => ENABLE, A => n175, ZN => n111);
   U46 : NAND2_X1 port map( A1 => D(20), A2 => ENABLE, ZN => n175);
   U47 : OAI21_X1 port map( B1 => n142, B2 => ENABLE, A => n174, ZN => n110);
   U48 : NAND2_X1 port map( A1 => D(21), A2 => ENABLE, ZN => n174);
   U49 : OAI21_X1 port map( B1 => n141, B2 => ENABLE, A => n173, ZN => n109);
   U50 : NAND2_X1 port map( A1 => D(22), A2 => ENABLE, ZN => n173);
   U51 : OAI21_X1 port map( B1 => n140, B2 => ENABLE, A => n172, ZN => n108);
   U52 : NAND2_X1 port map( A1 => D(23), A2 => ENABLE, ZN => n172);
   U53 : OAI21_X1 port map( B1 => n139, B2 => ENABLE, A => n171, ZN => n107);
   U54 : NAND2_X1 port map( A1 => D(24), A2 => ENABLE, ZN => n171);
   U55 : OAI21_X1 port map( B1 => n138, B2 => ENABLE, A => n170, ZN => n106);
   U56 : NAND2_X1 port map( A1 => D(25), A2 => ENABLE, ZN => n170);
   U57 : OAI21_X1 port map( B1 => n137, B2 => ENABLE, A => n169, ZN => n105);
   U58 : NAND2_X1 port map( A1 => D(26), A2 => ENABLE, ZN => n169);
   U59 : OAI21_X1 port map( B1 => n136, B2 => ENABLE, A => n168, ZN => n104);
   U60 : NAND2_X1 port map( A1 => D(27), A2 => ENABLE, ZN => n168);
   U61 : OAI21_X1 port map( B1 => n135, B2 => ENABLE, A => n167, ZN => n103);
   U62 : NAND2_X1 port map( A1 => D(28), A2 => ENABLE, ZN => n167);
   U63 : OAI21_X1 port map( B1 => n134, B2 => ENABLE, A => n166, ZN => n102);
   U64 : NAND2_X1 port map( A1 => D(29), A2 => ENABLE, ZN => n166);
   U65 : OAI21_X1 port map( B1 => n133, B2 => ENABLE, A => n165, ZN => n101);
   U66 : NAND2_X1 port map( A1 => D(30), A2 => ENABLE, ZN => n165);
   U67 : OAI21_X1 port map( B1 => n132, B2 => ENABLE, A => n164, ZN => n100);
   U68 : NAND2_X1 port map( A1 => D(31), A2 => ENABLE, ZN => n164);

end SYN_ASYNCHBEHAV;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity regFFD_NBIT32_11 is

   port( CK, RESET, ENABLE : in std_logic;  D : in std_logic_vector (31 downto 
         0);  Q : out std_logic_vector (31 downto 0));

end regFFD_NBIT32_11;

architecture SYN_ASYNCHBEHAV of regFFD_NBIT32_11 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, 
      n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, 
      n121, n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, 
      n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, 
      n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, 
      n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, 
      n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, 
      n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, 
      n193, n194, n195 : std_logic;

begin
   
   Q_reg_31_inst : DFFR_X1 port map( D => n100, CK => CK, RN => n99, Q => Q(31)
                           , QN => n132);
   Q_reg_30_inst : DFFR_X1 port map( D => n101, CK => CK, RN => n99, Q => Q(30)
                           , QN => n133);
   Q_reg_29_inst : DFFR_X1 port map( D => n102, CK => CK, RN => n99, Q => Q(29)
                           , QN => n134);
   Q_reg_28_inst : DFFR_X1 port map( D => n103, CK => CK, RN => n99, Q => Q(28)
                           , QN => n135);
   Q_reg_27_inst : DFFR_X1 port map( D => n104, CK => CK, RN => n99, Q => Q(27)
                           , QN => n136);
   Q_reg_26_inst : DFFR_X1 port map( D => n105, CK => CK, RN => n99, Q => Q(26)
                           , QN => n137);
   Q_reg_25_inst : DFFR_X1 port map( D => n106, CK => CK, RN => n99, Q => Q(25)
                           , QN => n138);
   Q_reg_24_inst : DFFR_X1 port map( D => n107, CK => CK, RN => n99, Q => Q(24)
                           , QN => n139);
   Q_reg_23_inst : DFFR_X1 port map( D => n108, CK => CK, RN => n98, Q => Q(23)
                           , QN => n140);
   Q_reg_22_inst : DFFR_X1 port map( D => n109, CK => CK, RN => n98, Q => Q(22)
                           , QN => n141);
   Q_reg_21_inst : DFFR_X1 port map( D => n110, CK => CK, RN => n98, Q => Q(21)
                           , QN => n142);
   Q_reg_20_inst : DFFR_X1 port map( D => n111, CK => CK, RN => n98, Q => Q(20)
                           , QN => n143);
   Q_reg_19_inst : DFFR_X1 port map( D => n112, CK => CK, RN => n98, Q => Q(19)
                           , QN => n144);
   Q_reg_18_inst : DFFR_X1 port map( D => n113, CK => CK, RN => n98, Q => Q(18)
                           , QN => n145);
   Q_reg_17_inst : DFFR_X1 port map( D => n114, CK => CK, RN => n98, Q => Q(17)
                           , QN => n146);
   Q_reg_16_inst : DFFR_X1 port map( D => n115, CK => CK, RN => n98, Q => Q(16)
                           , QN => n147);
   Q_reg_15_inst : DFFR_X1 port map( D => n116, CK => CK, RN => n98, Q => Q(15)
                           , QN => n148);
   Q_reg_14_inst : DFFR_X1 port map( D => n117, CK => CK, RN => n98, Q => Q(14)
                           , QN => n149);
   Q_reg_13_inst : DFFR_X1 port map( D => n118, CK => CK, RN => n98, Q => Q(13)
                           , QN => n150);
   Q_reg_12_inst : DFFR_X1 port map( D => n119, CK => CK, RN => n98, Q => Q(12)
                           , QN => n151);
   Q_reg_11_inst : DFFR_X1 port map( D => n120, CK => CK, RN => n97, Q => Q(11)
                           , QN => n152);
   Q_reg_10_inst : DFFR_X1 port map( D => n121, CK => CK, RN => n97, Q => Q(10)
                           , QN => n153);
   Q_reg_9_inst : DFFR_X1 port map( D => n122, CK => CK, RN => n97, Q => Q(9), 
                           QN => n154);
   Q_reg_8_inst : DFFR_X1 port map( D => n123, CK => CK, RN => n97, Q => Q(8), 
                           QN => n155);
   Q_reg_7_inst : DFFR_X1 port map( D => n124, CK => CK, RN => n97, Q => Q(7), 
                           QN => n156);
   Q_reg_6_inst : DFFR_X1 port map( D => n125, CK => CK, RN => n97, Q => Q(6), 
                           QN => n157);
   Q_reg_5_inst : DFFR_X1 port map( D => n126, CK => CK, RN => n97, Q => Q(5), 
                           QN => n158);
   Q_reg_4_inst : DFFR_X1 port map( D => n127, CK => CK, RN => n97, Q => Q(4), 
                           QN => n159);
   Q_reg_3_inst : DFFR_X1 port map( D => n128, CK => CK, RN => n97, Q => Q(3), 
                           QN => n160);
   Q_reg_2_inst : DFFR_X1 port map( D => n129, CK => CK, RN => n97, Q => Q(2), 
                           QN => n161);
   Q_reg_1_inst : DFFR_X1 port map( D => n130, CK => CK, RN => n97, Q => Q(1), 
                           QN => n162);
   Q_reg_0_inst : DFFR_X1 port map( D => n131, CK => CK, RN => n97, Q => Q(0), 
                           QN => n163);
   U2 : BUF_X1 port map( A => RESET, Z => n97);
   U3 : BUF_X1 port map( A => RESET, Z => n98);
   U4 : BUF_X1 port map( A => RESET, Z => n99);
   U5 : OAI21_X1 port map( B1 => n163, B2 => ENABLE, A => n195, ZN => n131);
   U6 : NAND2_X1 port map( A1 => ENABLE, A2 => D(0), ZN => n195);
   U7 : OAI21_X1 port map( B1 => n162, B2 => ENABLE, A => n194, ZN => n130);
   U8 : NAND2_X1 port map( A1 => D(1), A2 => ENABLE, ZN => n194);
   U9 : OAI21_X1 port map( B1 => n161, B2 => ENABLE, A => n193, ZN => n129);
   U10 : NAND2_X1 port map( A1 => D(2), A2 => ENABLE, ZN => n193);
   U11 : OAI21_X1 port map( B1 => n160, B2 => ENABLE, A => n192, ZN => n128);
   U12 : NAND2_X1 port map( A1 => D(3), A2 => ENABLE, ZN => n192);
   U13 : OAI21_X1 port map( B1 => n159, B2 => ENABLE, A => n191, ZN => n127);
   U14 : NAND2_X1 port map( A1 => D(4), A2 => ENABLE, ZN => n191);
   U15 : OAI21_X1 port map( B1 => n158, B2 => ENABLE, A => n190, ZN => n126);
   U16 : NAND2_X1 port map( A1 => D(5), A2 => ENABLE, ZN => n190);
   U17 : OAI21_X1 port map( B1 => n157, B2 => ENABLE, A => n189, ZN => n125);
   U18 : NAND2_X1 port map( A1 => D(6), A2 => ENABLE, ZN => n189);
   U19 : OAI21_X1 port map( B1 => n156, B2 => ENABLE, A => n188, ZN => n124);
   U20 : NAND2_X1 port map( A1 => D(7), A2 => ENABLE, ZN => n188);
   U21 : OAI21_X1 port map( B1 => n155, B2 => ENABLE, A => n187, ZN => n123);
   U22 : NAND2_X1 port map( A1 => D(8), A2 => ENABLE, ZN => n187);
   U23 : OAI21_X1 port map( B1 => n154, B2 => ENABLE, A => n186, ZN => n122);
   U24 : NAND2_X1 port map( A1 => D(9), A2 => ENABLE, ZN => n186);
   U25 : OAI21_X1 port map( B1 => n153, B2 => ENABLE, A => n185, ZN => n121);
   U26 : NAND2_X1 port map( A1 => D(10), A2 => ENABLE, ZN => n185);
   U27 : OAI21_X1 port map( B1 => n152, B2 => ENABLE, A => n184, ZN => n120);
   U28 : NAND2_X1 port map( A1 => D(11), A2 => ENABLE, ZN => n184);
   U29 : OAI21_X1 port map( B1 => n151, B2 => ENABLE, A => n183, ZN => n119);
   U30 : NAND2_X1 port map( A1 => D(12), A2 => ENABLE, ZN => n183);
   U31 : OAI21_X1 port map( B1 => n150, B2 => ENABLE, A => n182, ZN => n118);
   U32 : NAND2_X1 port map( A1 => D(13), A2 => ENABLE, ZN => n182);
   U33 : OAI21_X1 port map( B1 => n149, B2 => ENABLE, A => n181, ZN => n117);
   U34 : NAND2_X1 port map( A1 => D(14), A2 => ENABLE, ZN => n181);
   U35 : OAI21_X1 port map( B1 => n148, B2 => ENABLE, A => n180, ZN => n116);
   U36 : NAND2_X1 port map( A1 => D(15), A2 => ENABLE, ZN => n180);
   U37 : OAI21_X1 port map( B1 => n147, B2 => ENABLE, A => n179, ZN => n115);
   U38 : NAND2_X1 port map( A1 => D(16), A2 => ENABLE, ZN => n179);
   U39 : OAI21_X1 port map( B1 => n146, B2 => ENABLE, A => n178, ZN => n114);
   U40 : NAND2_X1 port map( A1 => D(17), A2 => ENABLE, ZN => n178);
   U41 : OAI21_X1 port map( B1 => n145, B2 => ENABLE, A => n177, ZN => n113);
   U42 : NAND2_X1 port map( A1 => D(18), A2 => ENABLE, ZN => n177);
   U43 : OAI21_X1 port map( B1 => n144, B2 => ENABLE, A => n176, ZN => n112);
   U44 : NAND2_X1 port map( A1 => D(19), A2 => ENABLE, ZN => n176);
   U45 : OAI21_X1 port map( B1 => n143, B2 => ENABLE, A => n175, ZN => n111);
   U46 : NAND2_X1 port map( A1 => D(20), A2 => ENABLE, ZN => n175);
   U47 : OAI21_X1 port map( B1 => n142, B2 => ENABLE, A => n174, ZN => n110);
   U48 : NAND2_X1 port map( A1 => D(21), A2 => ENABLE, ZN => n174);
   U49 : OAI21_X1 port map( B1 => n141, B2 => ENABLE, A => n173, ZN => n109);
   U50 : NAND2_X1 port map( A1 => D(22), A2 => ENABLE, ZN => n173);
   U51 : OAI21_X1 port map( B1 => n140, B2 => ENABLE, A => n172, ZN => n108);
   U52 : NAND2_X1 port map( A1 => D(23), A2 => ENABLE, ZN => n172);
   U53 : OAI21_X1 port map( B1 => n139, B2 => ENABLE, A => n171, ZN => n107);
   U54 : NAND2_X1 port map( A1 => D(24), A2 => ENABLE, ZN => n171);
   U55 : OAI21_X1 port map( B1 => n138, B2 => ENABLE, A => n170, ZN => n106);
   U56 : NAND2_X1 port map( A1 => D(25), A2 => ENABLE, ZN => n170);
   U57 : OAI21_X1 port map( B1 => n137, B2 => ENABLE, A => n169, ZN => n105);
   U58 : NAND2_X1 port map( A1 => D(26), A2 => ENABLE, ZN => n169);
   U59 : OAI21_X1 port map( B1 => n136, B2 => ENABLE, A => n168, ZN => n104);
   U60 : NAND2_X1 port map( A1 => D(27), A2 => ENABLE, ZN => n168);
   U61 : OAI21_X1 port map( B1 => n135, B2 => ENABLE, A => n167, ZN => n103);
   U62 : NAND2_X1 port map( A1 => D(28), A2 => ENABLE, ZN => n167);
   U63 : OAI21_X1 port map( B1 => n134, B2 => ENABLE, A => n166, ZN => n102);
   U64 : NAND2_X1 port map( A1 => D(29), A2 => ENABLE, ZN => n166);
   U65 : OAI21_X1 port map( B1 => n133, B2 => ENABLE, A => n165, ZN => n101);
   U66 : NAND2_X1 port map( A1 => D(30), A2 => ENABLE, ZN => n165);
   U67 : OAI21_X1 port map( B1 => n132, B2 => ENABLE, A => n164, ZN => n100);
   U68 : NAND2_X1 port map( A1 => D(31), A2 => ENABLE, ZN => n164);

end SYN_ASYNCHBEHAV;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity regFFD_NBIT32_10 is

   port( CK, RESET, ENABLE : in std_logic;  D : in std_logic_vector (31 downto 
         0);  Q : out std_logic_vector (31 downto 0));

end regFFD_NBIT32_10;

architecture SYN_ASYNCHBEHAV of regFFD_NBIT32_10 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, 
      n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, 
      n121, n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, 
      n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, 
      n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, 
      n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, 
      n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, 
      n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, 
      n193, n194, n195 : std_logic;

begin
   
   Q_reg_31_inst : DFFR_X1 port map( D => n100, CK => CK, RN => n99, Q => Q(31)
                           , QN => n132);
   Q_reg_30_inst : DFFR_X1 port map( D => n101, CK => CK, RN => n99, Q => Q(30)
                           , QN => n133);
   Q_reg_29_inst : DFFR_X1 port map( D => n102, CK => CK, RN => n99, Q => Q(29)
                           , QN => n134);
   Q_reg_28_inst : DFFR_X1 port map( D => n103, CK => CK, RN => n99, Q => Q(28)
                           , QN => n135);
   Q_reg_27_inst : DFFR_X1 port map( D => n104, CK => CK, RN => n99, Q => Q(27)
                           , QN => n136);
   Q_reg_26_inst : DFFR_X1 port map( D => n105, CK => CK, RN => n99, Q => Q(26)
                           , QN => n137);
   Q_reg_25_inst : DFFR_X1 port map( D => n106, CK => CK, RN => n99, Q => Q(25)
                           , QN => n138);
   Q_reg_24_inst : DFFR_X1 port map( D => n107, CK => CK, RN => n99, Q => Q(24)
                           , QN => n139);
   Q_reg_23_inst : DFFR_X1 port map( D => n108, CK => CK, RN => n98, Q => Q(23)
                           , QN => n140);
   Q_reg_22_inst : DFFR_X1 port map( D => n109, CK => CK, RN => n98, Q => Q(22)
                           , QN => n141);
   Q_reg_21_inst : DFFR_X1 port map( D => n110, CK => CK, RN => n98, Q => Q(21)
                           , QN => n142);
   Q_reg_20_inst : DFFR_X1 port map( D => n111, CK => CK, RN => n98, Q => Q(20)
                           , QN => n143);
   Q_reg_19_inst : DFFR_X1 port map( D => n112, CK => CK, RN => n98, Q => Q(19)
                           , QN => n144);
   Q_reg_18_inst : DFFR_X1 port map( D => n113, CK => CK, RN => n98, Q => Q(18)
                           , QN => n145);
   Q_reg_17_inst : DFFR_X1 port map( D => n114, CK => CK, RN => n98, Q => Q(17)
                           , QN => n146);
   Q_reg_16_inst : DFFR_X1 port map( D => n115, CK => CK, RN => n98, Q => Q(16)
                           , QN => n147);
   Q_reg_15_inst : DFFR_X1 port map( D => n116, CK => CK, RN => n98, Q => Q(15)
                           , QN => n148);
   Q_reg_14_inst : DFFR_X1 port map( D => n117, CK => CK, RN => n98, Q => Q(14)
                           , QN => n149);
   Q_reg_13_inst : DFFR_X1 port map( D => n118, CK => CK, RN => n98, Q => Q(13)
                           , QN => n150);
   Q_reg_12_inst : DFFR_X1 port map( D => n119, CK => CK, RN => n98, Q => Q(12)
                           , QN => n151);
   Q_reg_11_inst : DFFR_X1 port map( D => n120, CK => CK, RN => n97, Q => Q(11)
                           , QN => n152);
   Q_reg_10_inst : DFFR_X1 port map( D => n121, CK => CK, RN => n97, Q => Q(10)
                           , QN => n153);
   Q_reg_9_inst : DFFR_X1 port map( D => n122, CK => CK, RN => n97, Q => Q(9), 
                           QN => n154);
   Q_reg_8_inst : DFFR_X1 port map( D => n123, CK => CK, RN => n97, Q => Q(8), 
                           QN => n155);
   Q_reg_7_inst : DFFR_X1 port map( D => n124, CK => CK, RN => n97, Q => Q(7), 
                           QN => n156);
   Q_reg_6_inst : DFFR_X1 port map( D => n125, CK => CK, RN => n97, Q => Q(6), 
                           QN => n157);
   Q_reg_5_inst : DFFR_X1 port map( D => n126, CK => CK, RN => n97, Q => Q(5), 
                           QN => n158);
   Q_reg_4_inst : DFFR_X1 port map( D => n127, CK => CK, RN => n97, Q => Q(4), 
                           QN => n159);
   Q_reg_3_inst : DFFR_X1 port map( D => n128, CK => CK, RN => n97, Q => Q(3), 
                           QN => n160);
   Q_reg_2_inst : DFFR_X1 port map( D => n129, CK => CK, RN => n97, Q => Q(2), 
                           QN => n161);
   Q_reg_1_inst : DFFR_X1 port map( D => n130, CK => CK, RN => n97, Q => Q(1), 
                           QN => n162);
   Q_reg_0_inst : DFFR_X1 port map( D => n131, CK => CK, RN => n97, Q => Q(0), 
                           QN => n163);
   U2 : BUF_X1 port map( A => RESET, Z => n97);
   U3 : BUF_X1 port map( A => RESET, Z => n98);
   U4 : BUF_X1 port map( A => RESET, Z => n99);
   U5 : OAI21_X1 port map( B1 => n163, B2 => ENABLE, A => n195, ZN => n131);
   U6 : NAND2_X1 port map( A1 => ENABLE, A2 => D(0), ZN => n195);
   U7 : OAI21_X1 port map( B1 => n162, B2 => ENABLE, A => n194, ZN => n130);
   U8 : NAND2_X1 port map( A1 => D(1), A2 => ENABLE, ZN => n194);
   U9 : OAI21_X1 port map( B1 => n161, B2 => ENABLE, A => n193, ZN => n129);
   U10 : NAND2_X1 port map( A1 => D(2), A2 => ENABLE, ZN => n193);
   U11 : OAI21_X1 port map( B1 => n160, B2 => ENABLE, A => n192, ZN => n128);
   U12 : NAND2_X1 port map( A1 => D(3), A2 => ENABLE, ZN => n192);
   U13 : OAI21_X1 port map( B1 => n159, B2 => ENABLE, A => n191, ZN => n127);
   U14 : NAND2_X1 port map( A1 => D(4), A2 => ENABLE, ZN => n191);
   U15 : OAI21_X1 port map( B1 => n158, B2 => ENABLE, A => n190, ZN => n126);
   U16 : NAND2_X1 port map( A1 => D(5), A2 => ENABLE, ZN => n190);
   U17 : OAI21_X1 port map( B1 => n157, B2 => ENABLE, A => n189, ZN => n125);
   U18 : NAND2_X1 port map( A1 => D(6), A2 => ENABLE, ZN => n189);
   U19 : OAI21_X1 port map( B1 => n156, B2 => ENABLE, A => n188, ZN => n124);
   U20 : NAND2_X1 port map( A1 => D(7), A2 => ENABLE, ZN => n188);
   U21 : OAI21_X1 port map( B1 => n155, B2 => ENABLE, A => n187, ZN => n123);
   U22 : NAND2_X1 port map( A1 => D(8), A2 => ENABLE, ZN => n187);
   U23 : OAI21_X1 port map( B1 => n154, B2 => ENABLE, A => n186, ZN => n122);
   U24 : NAND2_X1 port map( A1 => D(9), A2 => ENABLE, ZN => n186);
   U25 : OAI21_X1 port map( B1 => n153, B2 => ENABLE, A => n185, ZN => n121);
   U26 : NAND2_X1 port map( A1 => D(10), A2 => ENABLE, ZN => n185);
   U27 : OAI21_X1 port map( B1 => n152, B2 => ENABLE, A => n184, ZN => n120);
   U28 : NAND2_X1 port map( A1 => D(11), A2 => ENABLE, ZN => n184);
   U29 : OAI21_X1 port map( B1 => n151, B2 => ENABLE, A => n183, ZN => n119);
   U30 : NAND2_X1 port map( A1 => D(12), A2 => ENABLE, ZN => n183);
   U31 : OAI21_X1 port map( B1 => n150, B2 => ENABLE, A => n182, ZN => n118);
   U32 : NAND2_X1 port map( A1 => D(13), A2 => ENABLE, ZN => n182);
   U33 : OAI21_X1 port map( B1 => n149, B2 => ENABLE, A => n181, ZN => n117);
   U34 : NAND2_X1 port map( A1 => D(14), A2 => ENABLE, ZN => n181);
   U35 : OAI21_X1 port map( B1 => n148, B2 => ENABLE, A => n180, ZN => n116);
   U36 : NAND2_X1 port map( A1 => D(15), A2 => ENABLE, ZN => n180);
   U37 : OAI21_X1 port map( B1 => n147, B2 => ENABLE, A => n179, ZN => n115);
   U38 : NAND2_X1 port map( A1 => D(16), A2 => ENABLE, ZN => n179);
   U39 : OAI21_X1 port map( B1 => n146, B2 => ENABLE, A => n178, ZN => n114);
   U40 : NAND2_X1 port map( A1 => D(17), A2 => ENABLE, ZN => n178);
   U41 : OAI21_X1 port map( B1 => n145, B2 => ENABLE, A => n177, ZN => n113);
   U42 : NAND2_X1 port map( A1 => D(18), A2 => ENABLE, ZN => n177);
   U43 : OAI21_X1 port map( B1 => n144, B2 => ENABLE, A => n176, ZN => n112);
   U44 : NAND2_X1 port map( A1 => D(19), A2 => ENABLE, ZN => n176);
   U45 : OAI21_X1 port map( B1 => n143, B2 => ENABLE, A => n175, ZN => n111);
   U46 : NAND2_X1 port map( A1 => D(20), A2 => ENABLE, ZN => n175);
   U47 : OAI21_X1 port map( B1 => n142, B2 => ENABLE, A => n174, ZN => n110);
   U48 : NAND2_X1 port map( A1 => D(21), A2 => ENABLE, ZN => n174);
   U49 : OAI21_X1 port map( B1 => n141, B2 => ENABLE, A => n173, ZN => n109);
   U50 : NAND2_X1 port map( A1 => D(22), A2 => ENABLE, ZN => n173);
   U51 : OAI21_X1 port map( B1 => n140, B2 => ENABLE, A => n172, ZN => n108);
   U52 : NAND2_X1 port map( A1 => D(23), A2 => ENABLE, ZN => n172);
   U53 : OAI21_X1 port map( B1 => n139, B2 => ENABLE, A => n171, ZN => n107);
   U54 : NAND2_X1 port map( A1 => D(24), A2 => ENABLE, ZN => n171);
   U55 : OAI21_X1 port map( B1 => n138, B2 => ENABLE, A => n170, ZN => n106);
   U56 : NAND2_X1 port map( A1 => D(25), A2 => ENABLE, ZN => n170);
   U57 : OAI21_X1 port map( B1 => n137, B2 => ENABLE, A => n169, ZN => n105);
   U58 : NAND2_X1 port map( A1 => D(26), A2 => ENABLE, ZN => n169);
   U59 : OAI21_X1 port map( B1 => n136, B2 => ENABLE, A => n168, ZN => n104);
   U60 : NAND2_X1 port map( A1 => D(27), A2 => ENABLE, ZN => n168);
   U61 : OAI21_X1 port map( B1 => n135, B2 => ENABLE, A => n167, ZN => n103);
   U62 : NAND2_X1 port map( A1 => D(28), A2 => ENABLE, ZN => n167);
   U63 : OAI21_X1 port map( B1 => n134, B2 => ENABLE, A => n166, ZN => n102);
   U64 : NAND2_X1 port map( A1 => D(29), A2 => ENABLE, ZN => n166);
   U65 : OAI21_X1 port map( B1 => n133, B2 => ENABLE, A => n165, ZN => n101);
   U66 : NAND2_X1 port map( A1 => D(30), A2 => ENABLE, ZN => n165);
   U67 : OAI21_X1 port map( B1 => n132, B2 => ENABLE, A => n164, ZN => n100);
   U68 : NAND2_X1 port map( A1 => D(31), A2 => ENABLE, ZN => n164);

end SYN_ASYNCHBEHAV;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity regFFD_NBIT32_9 is

   port( CK, RESET, ENABLE : in std_logic;  D : in std_logic_vector (31 downto 
         0);  Q : out std_logic_vector (31 downto 0));

end regFFD_NBIT32_9;

architecture SYN_ASYNCHBEHAV of regFFD_NBIT32_9 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, 
      n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, 
      n121, n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, 
      n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, 
      n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, 
      n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, 
      n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, 
      n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, 
      n193, n194, n195 : std_logic;

begin
   
   Q_reg_31_inst : DFFR_X1 port map( D => n100, CK => CK, RN => n99, Q => Q(31)
                           , QN => n132);
   Q_reg_30_inst : DFFR_X1 port map( D => n101, CK => CK, RN => n99, Q => Q(30)
                           , QN => n133);
   Q_reg_29_inst : DFFR_X1 port map( D => n102, CK => CK, RN => n99, Q => Q(29)
                           , QN => n134);
   Q_reg_28_inst : DFFR_X1 port map( D => n103, CK => CK, RN => n99, Q => Q(28)
                           , QN => n135);
   Q_reg_27_inst : DFFR_X1 port map( D => n104, CK => CK, RN => n99, Q => Q(27)
                           , QN => n136);
   Q_reg_26_inst : DFFR_X1 port map( D => n105, CK => CK, RN => n99, Q => Q(26)
                           , QN => n137);
   Q_reg_25_inst : DFFR_X1 port map( D => n106, CK => CK, RN => n99, Q => Q(25)
                           , QN => n138);
   Q_reg_24_inst : DFFR_X1 port map( D => n107, CK => CK, RN => n99, Q => Q(24)
                           , QN => n139);
   Q_reg_23_inst : DFFR_X1 port map( D => n108, CK => CK, RN => n98, Q => Q(23)
                           , QN => n140);
   Q_reg_22_inst : DFFR_X1 port map( D => n109, CK => CK, RN => n98, Q => Q(22)
                           , QN => n141);
   Q_reg_21_inst : DFFR_X1 port map( D => n110, CK => CK, RN => n98, Q => Q(21)
                           , QN => n142);
   Q_reg_20_inst : DFFR_X1 port map( D => n111, CK => CK, RN => n98, Q => Q(20)
                           , QN => n143);
   Q_reg_19_inst : DFFR_X1 port map( D => n112, CK => CK, RN => n98, Q => Q(19)
                           , QN => n144);
   Q_reg_18_inst : DFFR_X1 port map( D => n113, CK => CK, RN => n98, Q => Q(18)
                           , QN => n145);
   Q_reg_17_inst : DFFR_X1 port map( D => n114, CK => CK, RN => n98, Q => Q(17)
                           , QN => n146);
   Q_reg_16_inst : DFFR_X1 port map( D => n115, CK => CK, RN => n98, Q => Q(16)
                           , QN => n147);
   Q_reg_15_inst : DFFR_X1 port map( D => n116, CK => CK, RN => n98, Q => Q(15)
                           , QN => n148);
   Q_reg_14_inst : DFFR_X1 port map( D => n117, CK => CK, RN => n98, Q => Q(14)
                           , QN => n149);
   Q_reg_13_inst : DFFR_X1 port map( D => n118, CK => CK, RN => n98, Q => Q(13)
                           , QN => n150);
   Q_reg_12_inst : DFFR_X1 port map( D => n119, CK => CK, RN => n98, Q => Q(12)
                           , QN => n151);
   Q_reg_11_inst : DFFR_X1 port map( D => n120, CK => CK, RN => n97, Q => Q(11)
                           , QN => n152);
   Q_reg_10_inst : DFFR_X1 port map( D => n121, CK => CK, RN => n97, Q => Q(10)
                           , QN => n153);
   Q_reg_9_inst : DFFR_X1 port map( D => n122, CK => CK, RN => n97, Q => Q(9), 
                           QN => n154);
   Q_reg_8_inst : DFFR_X1 port map( D => n123, CK => CK, RN => n97, Q => Q(8), 
                           QN => n155);
   Q_reg_7_inst : DFFR_X1 port map( D => n124, CK => CK, RN => n97, Q => Q(7), 
                           QN => n156);
   Q_reg_6_inst : DFFR_X1 port map( D => n125, CK => CK, RN => n97, Q => Q(6), 
                           QN => n157);
   Q_reg_5_inst : DFFR_X1 port map( D => n126, CK => CK, RN => n97, Q => Q(5), 
                           QN => n158);
   Q_reg_4_inst : DFFR_X1 port map( D => n127, CK => CK, RN => n97, Q => Q(4), 
                           QN => n159);
   Q_reg_3_inst : DFFR_X1 port map( D => n128, CK => CK, RN => n97, Q => Q(3), 
                           QN => n160);
   Q_reg_2_inst : DFFR_X1 port map( D => n129, CK => CK, RN => n97, Q => Q(2), 
                           QN => n161);
   Q_reg_1_inst : DFFR_X1 port map( D => n130, CK => CK, RN => n97, Q => Q(1), 
                           QN => n162);
   Q_reg_0_inst : DFFR_X1 port map( D => n131, CK => CK, RN => n97, Q => Q(0), 
                           QN => n163);
   U2 : BUF_X1 port map( A => RESET, Z => n97);
   U3 : BUF_X1 port map( A => RESET, Z => n98);
   U4 : BUF_X1 port map( A => RESET, Z => n99);
   U5 : OAI21_X1 port map( B1 => n163, B2 => ENABLE, A => n195, ZN => n131);
   U6 : NAND2_X1 port map( A1 => ENABLE, A2 => D(0), ZN => n195);
   U7 : OAI21_X1 port map( B1 => n162, B2 => ENABLE, A => n194, ZN => n130);
   U8 : NAND2_X1 port map( A1 => D(1), A2 => ENABLE, ZN => n194);
   U9 : OAI21_X1 port map( B1 => n161, B2 => ENABLE, A => n193, ZN => n129);
   U10 : NAND2_X1 port map( A1 => D(2), A2 => ENABLE, ZN => n193);
   U11 : OAI21_X1 port map( B1 => n160, B2 => ENABLE, A => n192, ZN => n128);
   U12 : NAND2_X1 port map( A1 => D(3), A2 => ENABLE, ZN => n192);
   U13 : OAI21_X1 port map( B1 => n159, B2 => ENABLE, A => n191, ZN => n127);
   U14 : NAND2_X1 port map( A1 => D(4), A2 => ENABLE, ZN => n191);
   U15 : OAI21_X1 port map( B1 => n158, B2 => ENABLE, A => n190, ZN => n126);
   U16 : NAND2_X1 port map( A1 => D(5), A2 => ENABLE, ZN => n190);
   U17 : OAI21_X1 port map( B1 => n157, B2 => ENABLE, A => n189, ZN => n125);
   U18 : NAND2_X1 port map( A1 => D(6), A2 => ENABLE, ZN => n189);
   U19 : OAI21_X1 port map( B1 => n156, B2 => ENABLE, A => n188, ZN => n124);
   U20 : NAND2_X1 port map( A1 => D(7), A2 => ENABLE, ZN => n188);
   U21 : OAI21_X1 port map( B1 => n155, B2 => ENABLE, A => n187, ZN => n123);
   U22 : NAND2_X1 port map( A1 => D(8), A2 => ENABLE, ZN => n187);
   U23 : OAI21_X1 port map( B1 => n154, B2 => ENABLE, A => n186, ZN => n122);
   U24 : NAND2_X1 port map( A1 => D(9), A2 => ENABLE, ZN => n186);
   U25 : OAI21_X1 port map( B1 => n153, B2 => ENABLE, A => n185, ZN => n121);
   U26 : NAND2_X1 port map( A1 => D(10), A2 => ENABLE, ZN => n185);
   U27 : OAI21_X1 port map( B1 => n152, B2 => ENABLE, A => n184, ZN => n120);
   U28 : NAND2_X1 port map( A1 => D(11), A2 => ENABLE, ZN => n184);
   U29 : OAI21_X1 port map( B1 => n151, B2 => ENABLE, A => n183, ZN => n119);
   U30 : NAND2_X1 port map( A1 => D(12), A2 => ENABLE, ZN => n183);
   U31 : OAI21_X1 port map( B1 => n150, B2 => ENABLE, A => n182, ZN => n118);
   U32 : NAND2_X1 port map( A1 => D(13), A2 => ENABLE, ZN => n182);
   U33 : OAI21_X1 port map( B1 => n149, B2 => ENABLE, A => n181, ZN => n117);
   U34 : NAND2_X1 port map( A1 => D(14), A2 => ENABLE, ZN => n181);
   U35 : OAI21_X1 port map( B1 => n148, B2 => ENABLE, A => n180, ZN => n116);
   U36 : NAND2_X1 port map( A1 => D(15), A2 => ENABLE, ZN => n180);
   U37 : OAI21_X1 port map( B1 => n147, B2 => ENABLE, A => n179, ZN => n115);
   U38 : NAND2_X1 port map( A1 => D(16), A2 => ENABLE, ZN => n179);
   U39 : OAI21_X1 port map( B1 => n146, B2 => ENABLE, A => n178, ZN => n114);
   U40 : NAND2_X1 port map( A1 => D(17), A2 => ENABLE, ZN => n178);
   U41 : OAI21_X1 port map( B1 => n145, B2 => ENABLE, A => n177, ZN => n113);
   U42 : NAND2_X1 port map( A1 => D(18), A2 => ENABLE, ZN => n177);
   U43 : OAI21_X1 port map( B1 => n144, B2 => ENABLE, A => n176, ZN => n112);
   U44 : NAND2_X1 port map( A1 => D(19), A2 => ENABLE, ZN => n176);
   U45 : OAI21_X1 port map( B1 => n143, B2 => ENABLE, A => n175, ZN => n111);
   U46 : NAND2_X1 port map( A1 => D(20), A2 => ENABLE, ZN => n175);
   U47 : OAI21_X1 port map( B1 => n142, B2 => ENABLE, A => n174, ZN => n110);
   U48 : NAND2_X1 port map( A1 => D(21), A2 => ENABLE, ZN => n174);
   U49 : OAI21_X1 port map( B1 => n141, B2 => ENABLE, A => n173, ZN => n109);
   U50 : NAND2_X1 port map( A1 => D(22), A2 => ENABLE, ZN => n173);
   U51 : OAI21_X1 port map( B1 => n140, B2 => ENABLE, A => n172, ZN => n108);
   U52 : NAND2_X1 port map( A1 => D(23), A2 => ENABLE, ZN => n172);
   U53 : OAI21_X1 port map( B1 => n139, B2 => ENABLE, A => n171, ZN => n107);
   U54 : NAND2_X1 port map( A1 => D(24), A2 => ENABLE, ZN => n171);
   U55 : OAI21_X1 port map( B1 => n138, B2 => ENABLE, A => n170, ZN => n106);
   U56 : NAND2_X1 port map( A1 => D(25), A2 => ENABLE, ZN => n170);
   U57 : OAI21_X1 port map( B1 => n137, B2 => ENABLE, A => n169, ZN => n105);
   U58 : NAND2_X1 port map( A1 => D(26), A2 => ENABLE, ZN => n169);
   U59 : OAI21_X1 port map( B1 => n136, B2 => ENABLE, A => n168, ZN => n104);
   U60 : NAND2_X1 port map( A1 => D(27), A2 => ENABLE, ZN => n168);
   U61 : OAI21_X1 port map( B1 => n135, B2 => ENABLE, A => n167, ZN => n103);
   U62 : NAND2_X1 port map( A1 => D(28), A2 => ENABLE, ZN => n167);
   U63 : OAI21_X1 port map( B1 => n134, B2 => ENABLE, A => n166, ZN => n102);
   U64 : NAND2_X1 port map( A1 => D(29), A2 => ENABLE, ZN => n166);
   U65 : OAI21_X1 port map( B1 => n133, B2 => ENABLE, A => n165, ZN => n101);
   U66 : NAND2_X1 port map( A1 => D(30), A2 => ENABLE, ZN => n165);
   U67 : OAI21_X1 port map( B1 => n132, B2 => ENABLE, A => n164, ZN => n100);
   U68 : NAND2_X1 port map( A1 => D(31), A2 => ENABLE, ZN => n164);

end SYN_ASYNCHBEHAV;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity regFFD_NBIT32_8 is

   port( CK, RESET, ENABLE : in std_logic;  D : in std_logic_vector (31 downto 
         0);  Q : out std_logic_vector (31 downto 0));

end regFFD_NBIT32_8;

architecture SYN_ASYNCHBEHAV of regFFD_NBIT32_8 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, 
      n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, 
      n121, n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, 
      n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, 
      n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, 
      n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, 
      n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, 
      n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, 
      n193, n194, n195 : std_logic;

begin
   
   Q_reg_31_inst : DFFR_X1 port map( D => n100, CK => CK, RN => n99, Q => Q(31)
                           , QN => n132);
   Q_reg_30_inst : DFFR_X1 port map( D => n101, CK => CK, RN => n99, Q => Q(30)
                           , QN => n133);
   Q_reg_29_inst : DFFR_X1 port map( D => n102, CK => CK, RN => n99, Q => Q(29)
                           , QN => n134);
   Q_reg_28_inst : DFFR_X1 port map( D => n103, CK => CK, RN => n99, Q => Q(28)
                           , QN => n135);
   Q_reg_27_inst : DFFR_X1 port map( D => n104, CK => CK, RN => n99, Q => Q(27)
                           , QN => n136);
   Q_reg_26_inst : DFFR_X1 port map( D => n105, CK => CK, RN => n99, Q => Q(26)
                           , QN => n137);
   Q_reg_25_inst : DFFR_X1 port map( D => n106, CK => CK, RN => n99, Q => Q(25)
                           , QN => n138);
   Q_reg_24_inst : DFFR_X1 port map( D => n107, CK => CK, RN => n99, Q => Q(24)
                           , QN => n139);
   Q_reg_23_inst : DFFR_X1 port map( D => n108, CK => CK, RN => n98, Q => Q(23)
                           , QN => n140);
   Q_reg_22_inst : DFFR_X1 port map( D => n109, CK => CK, RN => n98, Q => Q(22)
                           , QN => n141);
   Q_reg_21_inst : DFFR_X1 port map( D => n110, CK => CK, RN => n98, Q => Q(21)
                           , QN => n142);
   Q_reg_20_inst : DFFR_X1 port map( D => n111, CK => CK, RN => n98, Q => Q(20)
                           , QN => n143);
   Q_reg_19_inst : DFFR_X1 port map( D => n112, CK => CK, RN => n98, Q => Q(19)
                           , QN => n144);
   Q_reg_18_inst : DFFR_X1 port map( D => n113, CK => CK, RN => n98, Q => Q(18)
                           , QN => n145);
   Q_reg_17_inst : DFFR_X1 port map( D => n114, CK => CK, RN => n98, Q => Q(17)
                           , QN => n146);
   Q_reg_16_inst : DFFR_X1 port map( D => n115, CK => CK, RN => n98, Q => Q(16)
                           , QN => n147);
   Q_reg_15_inst : DFFR_X1 port map( D => n116, CK => CK, RN => n98, Q => Q(15)
                           , QN => n148);
   Q_reg_14_inst : DFFR_X1 port map( D => n117, CK => CK, RN => n98, Q => Q(14)
                           , QN => n149);
   Q_reg_13_inst : DFFR_X1 port map( D => n118, CK => CK, RN => n98, Q => Q(13)
                           , QN => n150);
   Q_reg_12_inst : DFFR_X1 port map( D => n119, CK => CK, RN => n98, Q => Q(12)
                           , QN => n151);
   Q_reg_11_inst : DFFR_X1 port map( D => n120, CK => CK, RN => n97, Q => Q(11)
                           , QN => n152);
   Q_reg_10_inst : DFFR_X1 port map( D => n121, CK => CK, RN => n97, Q => Q(10)
                           , QN => n153);
   Q_reg_9_inst : DFFR_X1 port map( D => n122, CK => CK, RN => n97, Q => Q(9), 
                           QN => n154);
   Q_reg_8_inst : DFFR_X1 port map( D => n123, CK => CK, RN => n97, Q => Q(8), 
                           QN => n155);
   Q_reg_7_inst : DFFR_X1 port map( D => n124, CK => CK, RN => n97, Q => Q(7), 
                           QN => n156);
   Q_reg_6_inst : DFFR_X1 port map( D => n125, CK => CK, RN => n97, Q => Q(6), 
                           QN => n157);
   Q_reg_5_inst : DFFR_X1 port map( D => n126, CK => CK, RN => n97, Q => Q(5), 
                           QN => n158);
   Q_reg_4_inst : DFFR_X1 port map( D => n127, CK => CK, RN => n97, Q => Q(4), 
                           QN => n159);
   Q_reg_3_inst : DFFR_X1 port map( D => n128, CK => CK, RN => n97, Q => Q(3), 
                           QN => n160);
   Q_reg_2_inst : DFFR_X1 port map( D => n129, CK => CK, RN => n97, Q => Q(2), 
                           QN => n161);
   Q_reg_1_inst : DFFR_X1 port map( D => n130, CK => CK, RN => n97, Q => Q(1), 
                           QN => n162);
   Q_reg_0_inst : DFFR_X1 port map( D => n131, CK => CK, RN => n97, Q => Q(0), 
                           QN => n163);
   U2 : BUF_X1 port map( A => RESET, Z => n97);
   U3 : BUF_X1 port map( A => RESET, Z => n98);
   U4 : BUF_X1 port map( A => RESET, Z => n99);
   U5 : OAI21_X1 port map( B1 => n163, B2 => ENABLE, A => n195, ZN => n131);
   U6 : NAND2_X1 port map( A1 => ENABLE, A2 => D(0), ZN => n195);
   U7 : OAI21_X1 port map( B1 => n162, B2 => ENABLE, A => n194, ZN => n130);
   U8 : NAND2_X1 port map( A1 => D(1), A2 => ENABLE, ZN => n194);
   U9 : OAI21_X1 port map( B1 => n161, B2 => ENABLE, A => n193, ZN => n129);
   U10 : NAND2_X1 port map( A1 => D(2), A2 => ENABLE, ZN => n193);
   U11 : OAI21_X1 port map( B1 => n160, B2 => ENABLE, A => n192, ZN => n128);
   U12 : NAND2_X1 port map( A1 => D(3), A2 => ENABLE, ZN => n192);
   U13 : OAI21_X1 port map( B1 => n159, B2 => ENABLE, A => n191, ZN => n127);
   U14 : NAND2_X1 port map( A1 => D(4), A2 => ENABLE, ZN => n191);
   U15 : OAI21_X1 port map( B1 => n158, B2 => ENABLE, A => n190, ZN => n126);
   U16 : NAND2_X1 port map( A1 => D(5), A2 => ENABLE, ZN => n190);
   U17 : OAI21_X1 port map( B1 => n157, B2 => ENABLE, A => n189, ZN => n125);
   U18 : NAND2_X1 port map( A1 => D(6), A2 => ENABLE, ZN => n189);
   U19 : OAI21_X1 port map( B1 => n156, B2 => ENABLE, A => n188, ZN => n124);
   U20 : NAND2_X1 port map( A1 => D(7), A2 => ENABLE, ZN => n188);
   U21 : OAI21_X1 port map( B1 => n155, B2 => ENABLE, A => n187, ZN => n123);
   U22 : NAND2_X1 port map( A1 => D(8), A2 => ENABLE, ZN => n187);
   U23 : OAI21_X1 port map( B1 => n154, B2 => ENABLE, A => n186, ZN => n122);
   U24 : NAND2_X1 port map( A1 => D(9), A2 => ENABLE, ZN => n186);
   U25 : OAI21_X1 port map( B1 => n153, B2 => ENABLE, A => n185, ZN => n121);
   U26 : NAND2_X1 port map( A1 => D(10), A2 => ENABLE, ZN => n185);
   U27 : OAI21_X1 port map( B1 => n152, B2 => ENABLE, A => n184, ZN => n120);
   U28 : NAND2_X1 port map( A1 => D(11), A2 => ENABLE, ZN => n184);
   U29 : OAI21_X1 port map( B1 => n151, B2 => ENABLE, A => n183, ZN => n119);
   U30 : NAND2_X1 port map( A1 => D(12), A2 => ENABLE, ZN => n183);
   U31 : OAI21_X1 port map( B1 => n150, B2 => ENABLE, A => n182, ZN => n118);
   U32 : NAND2_X1 port map( A1 => D(13), A2 => ENABLE, ZN => n182);
   U33 : OAI21_X1 port map( B1 => n149, B2 => ENABLE, A => n181, ZN => n117);
   U34 : NAND2_X1 port map( A1 => D(14), A2 => ENABLE, ZN => n181);
   U35 : OAI21_X1 port map( B1 => n148, B2 => ENABLE, A => n180, ZN => n116);
   U36 : NAND2_X1 port map( A1 => D(15), A2 => ENABLE, ZN => n180);
   U37 : OAI21_X1 port map( B1 => n147, B2 => ENABLE, A => n179, ZN => n115);
   U38 : NAND2_X1 port map( A1 => D(16), A2 => ENABLE, ZN => n179);
   U39 : OAI21_X1 port map( B1 => n146, B2 => ENABLE, A => n178, ZN => n114);
   U40 : NAND2_X1 port map( A1 => D(17), A2 => ENABLE, ZN => n178);
   U41 : OAI21_X1 port map( B1 => n145, B2 => ENABLE, A => n177, ZN => n113);
   U42 : NAND2_X1 port map( A1 => D(18), A2 => ENABLE, ZN => n177);
   U43 : OAI21_X1 port map( B1 => n144, B2 => ENABLE, A => n176, ZN => n112);
   U44 : NAND2_X1 port map( A1 => D(19), A2 => ENABLE, ZN => n176);
   U45 : OAI21_X1 port map( B1 => n143, B2 => ENABLE, A => n175, ZN => n111);
   U46 : NAND2_X1 port map( A1 => D(20), A2 => ENABLE, ZN => n175);
   U47 : OAI21_X1 port map( B1 => n142, B2 => ENABLE, A => n174, ZN => n110);
   U48 : NAND2_X1 port map( A1 => D(21), A2 => ENABLE, ZN => n174);
   U49 : OAI21_X1 port map( B1 => n141, B2 => ENABLE, A => n173, ZN => n109);
   U50 : NAND2_X1 port map( A1 => D(22), A2 => ENABLE, ZN => n173);
   U51 : OAI21_X1 port map( B1 => n140, B2 => ENABLE, A => n172, ZN => n108);
   U52 : NAND2_X1 port map( A1 => D(23), A2 => ENABLE, ZN => n172);
   U53 : OAI21_X1 port map( B1 => n139, B2 => ENABLE, A => n171, ZN => n107);
   U54 : NAND2_X1 port map( A1 => D(24), A2 => ENABLE, ZN => n171);
   U55 : OAI21_X1 port map( B1 => n138, B2 => ENABLE, A => n170, ZN => n106);
   U56 : NAND2_X1 port map( A1 => D(25), A2 => ENABLE, ZN => n170);
   U57 : OAI21_X1 port map( B1 => n137, B2 => ENABLE, A => n169, ZN => n105);
   U58 : NAND2_X1 port map( A1 => D(26), A2 => ENABLE, ZN => n169);
   U59 : OAI21_X1 port map( B1 => n136, B2 => ENABLE, A => n168, ZN => n104);
   U60 : NAND2_X1 port map( A1 => D(27), A2 => ENABLE, ZN => n168);
   U61 : OAI21_X1 port map( B1 => n135, B2 => ENABLE, A => n167, ZN => n103);
   U62 : NAND2_X1 port map( A1 => D(28), A2 => ENABLE, ZN => n167);
   U63 : OAI21_X1 port map( B1 => n134, B2 => ENABLE, A => n166, ZN => n102);
   U64 : NAND2_X1 port map( A1 => D(29), A2 => ENABLE, ZN => n166);
   U65 : OAI21_X1 port map( B1 => n133, B2 => ENABLE, A => n165, ZN => n101);
   U66 : NAND2_X1 port map( A1 => D(30), A2 => ENABLE, ZN => n165);
   U67 : OAI21_X1 port map( B1 => n132, B2 => ENABLE, A => n164, ZN => n100);
   U68 : NAND2_X1 port map( A1 => D(31), A2 => ENABLE, ZN => n164);

end SYN_ASYNCHBEHAV;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity regFFD_NBIT32_7 is

   port( CK, RESET, ENABLE : in std_logic;  D : in std_logic_vector (31 downto 
         0);  Q : out std_logic_vector (31 downto 0));

end regFFD_NBIT32_7;

architecture SYN_ASYNCHBEHAV of regFFD_NBIT32_7 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, 
      n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, 
      n121, n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, 
      n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, 
      n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, 
      n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, 
      n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, 
      n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, 
      n193, n194, n195 : std_logic;

begin
   
   Q_reg_31_inst : DFFR_X1 port map( D => n100, CK => CK, RN => n99, Q => Q(31)
                           , QN => n132);
   Q_reg_30_inst : DFFR_X1 port map( D => n101, CK => CK, RN => n99, Q => Q(30)
                           , QN => n133);
   Q_reg_29_inst : DFFR_X1 port map( D => n102, CK => CK, RN => n99, Q => Q(29)
                           , QN => n134);
   Q_reg_28_inst : DFFR_X1 port map( D => n103, CK => CK, RN => n99, Q => Q(28)
                           , QN => n135);
   Q_reg_27_inst : DFFR_X1 port map( D => n104, CK => CK, RN => n99, Q => Q(27)
                           , QN => n136);
   Q_reg_26_inst : DFFR_X1 port map( D => n105, CK => CK, RN => n99, Q => Q(26)
                           , QN => n137);
   Q_reg_25_inst : DFFR_X1 port map( D => n106, CK => CK, RN => n99, Q => Q(25)
                           , QN => n138);
   Q_reg_24_inst : DFFR_X1 port map( D => n107, CK => CK, RN => n99, Q => Q(24)
                           , QN => n139);
   Q_reg_23_inst : DFFR_X1 port map( D => n108, CK => CK, RN => n98, Q => Q(23)
                           , QN => n140);
   Q_reg_22_inst : DFFR_X1 port map( D => n109, CK => CK, RN => n98, Q => Q(22)
                           , QN => n141);
   Q_reg_21_inst : DFFR_X1 port map( D => n110, CK => CK, RN => n98, Q => Q(21)
                           , QN => n142);
   Q_reg_20_inst : DFFR_X1 port map( D => n111, CK => CK, RN => n98, Q => Q(20)
                           , QN => n143);
   Q_reg_19_inst : DFFR_X1 port map( D => n112, CK => CK, RN => n98, Q => Q(19)
                           , QN => n144);
   Q_reg_18_inst : DFFR_X1 port map( D => n113, CK => CK, RN => n98, Q => Q(18)
                           , QN => n145);
   Q_reg_17_inst : DFFR_X1 port map( D => n114, CK => CK, RN => n98, Q => Q(17)
                           , QN => n146);
   Q_reg_16_inst : DFFR_X1 port map( D => n115, CK => CK, RN => n98, Q => Q(16)
                           , QN => n147);
   Q_reg_15_inst : DFFR_X1 port map( D => n116, CK => CK, RN => n98, Q => Q(15)
                           , QN => n148);
   Q_reg_14_inst : DFFR_X1 port map( D => n117, CK => CK, RN => n98, Q => Q(14)
                           , QN => n149);
   Q_reg_13_inst : DFFR_X1 port map( D => n118, CK => CK, RN => n98, Q => Q(13)
                           , QN => n150);
   Q_reg_12_inst : DFFR_X1 port map( D => n119, CK => CK, RN => n98, Q => Q(12)
                           , QN => n151);
   Q_reg_11_inst : DFFR_X1 port map( D => n120, CK => CK, RN => n97, Q => Q(11)
                           , QN => n152);
   Q_reg_10_inst : DFFR_X1 port map( D => n121, CK => CK, RN => n97, Q => Q(10)
                           , QN => n153);
   Q_reg_9_inst : DFFR_X1 port map( D => n122, CK => CK, RN => n97, Q => Q(9), 
                           QN => n154);
   Q_reg_8_inst : DFFR_X1 port map( D => n123, CK => CK, RN => n97, Q => Q(8), 
                           QN => n155);
   Q_reg_7_inst : DFFR_X1 port map( D => n124, CK => CK, RN => n97, Q => Q(7), 
                           QN => n156);
   Q_reg_6_inst : DFFR_X1 port map( D => n125, CK => CK, RN => n97, Q => Q(6), 
                           QN => n157);
   Q_reg_5_inst : DFFR_X1 port map( D => n126, CK => CK, RN => n97, Q => Q(5), 
                           QN => n158);
   Q_reg_4_inst : DFFR_X1 port map( D => n127, CK => CK, RN => n97, Q => Q(4), 
                           QN => n159);
   Q_reg_3_inst : DFFR_X1 port map( D => n128, CK => CK, RN => n97, Q => Q(3), 
                           QN => n160);
   Q_reg_2_inst : DFFR_X1 port map( D => n129, CK => CK, RN => n97, Q => Q(2), 
                           QN => n161);
   Q_reg_1_inst : DFFR_X1 port map( D => n130, CK => CK, RN => n97, Q => Q(1), 
                           QN => n162);
   Q_reg_0_inst : DFFR_X1 port map( D => n131, CK => CK, RN => n97, Q => Q(0), 
                           QN => n163);
   U2 : BUF_X1 port map( A => RESET, Z => n97);
   U3 : BUF_X1 port map( A => RESET, Z => n98);
   U4 : BUF_X1 port map( A => RESET, Z => n99);
   U5 : OAI21_X1 port map( B1 => n163, B2 => ENABLE, A => n195, ZN => n131);
   U6 : NAND2_X1 port map( A1 => ENABLE, A2 => D(0), ZN => n195);
   U7 : OAI21_X1 port map( B1 => n162, B2 => ENABLE, A => n194, ZN => n130);
   U8 : NAND2_X1 port map( A1 => D(1), A2 => ENABLE, ZN => n194);
   U9 : OAI21_X1 port map( B1 => n161, B2 => ENABLE, A => n193, ZN => n129);
   U10 : NAND2_X1 port map( A1 => D(2), A2 => ENABLE, ZN => n193);
   U11 : OAI21_X1 port map( B1 => n160, B2 => ENABLE, A => n192, ZN => n128);
   U12 : NAND2_X1 port map( A1 => D(3), A2 => ENABLE, ZN => n192);
   U13 : OAI21_X1 port map( B1 => n159, B2 => ENABLE, A => n191, ZN => n127);
   U14 : NAND2_X1 port map( A1 => D(4), A2 => ENABLE, ZN => n191);
   U15 : OAI21_X1 port map( B1 => n158, B2 => ENABLE, A => n190, ZN => n126);
   U16 : NAND2_X1 port map( A1 => D(5), A2 => ENABLE, ZN => n190);
   U17 : OAI21_X1 port map( B1 => n157, B2 => ENABLE, A => n189, ZN => n125);
   U18 : NAND2_X1 port map( A1 => D(6), A2 => ENABLE, ZN => n189);
   U19 : OAI21_X1 port map( B1 => n156, B2 => ENABLE, A => n188, ZN => n124);
   U20 : NAND2_X1 port map( A1 => D(7), A2 => ENABLE, ZN => n188);
   U21 : OAI21_X1 port map( B1 => n155, B2 => ENABLE, A => n187, ZN => n123);
   U22 : NAND2_X1 port map( A1 => D(8), A2 => ENABLE, ZN => n187);
   U23 : OAI21_X1 port map( B1 => n154, B2 => ENABLE, A => n186, ZN => n122);
   U24 : NAND2_X1 port map( A1 => D(9), A2 => ENABLE, ZN => n186);
   U25 : OAI21_X1 port map( B1 => n153, B2 => ENABLE, A => n185, ZN => n121);
   U26 : NAND2_X1 port map( A1 => D(10), A2 => ENABLE, ZN => n185);
   U27 : OAI21_X1 port map( B1 => n152, B2 => ENABLE, A => n184, ZN => n120);
   U28 : NAND2_X1 port map( A1 => D(11), A2 => ENABLE, ZN => n184);
   U29 : OAI21_X1 port map( B1 => n151, B2 => ENABLE, A => n183, ZN => n119);
   U30 : NAND2_X1 port map( A1 => D(12), A2 => ENABLE, ZN => n183);
   U31 : OAI21_X1 port map( B1 => n150, B2 => ENABLE, A => n182, ZN => n118);
   U32 : NAND2_X1 port map( A1 => D(13), A2 => ENABLE, ZN => n182);
   U33 : OAI21_X1 port map( B1 => n149, B2 => ENABLE, A => n181, ZN => n117);
   U34 : NAND2_X1 port map( A1 => D(14), A2 => ENABLE, ZN => n181);
   U35 : OAI21_X1 port map( B1 => n148, B2 => ENABLE, A => n180, ZN => n116);
   U36 : NAND2_X1 port map( A1 => D(15), A2 => ENABLE, ZN => n180);
   U37 : OAI21_X1 port map( B1 => n147, B2 => ENABLE, A => n179, ZN => n115);
   U38 : NAND2_X1 port map( A1 => D(16), A2 => ENABLE, ZN => n179);
   U39 : OAI21_X1 port map( B1 => n146, B2 => ENABLE, A => n178, ZN => n114);
   U40 : NAND2_X1 port map( A1 => D(17), A2 => ENABLE, ZN => n178);
   U41 : OAI21_X1 port map( B1 => n145, B2 => ENABLE, A => n177, ZN => n113);
   U42 : NAND2_X1 port map( A1 => D(18), A2 => ENABLE, ZN => n177);
   U43 : OAI21_X1 port map( B1 => n144, B2 => ENABLE, A => n176, ZN => n112);
   U44 : NAND2_X1 port map( A1 => D(19), A2 => ENABLE, ZN => n176);
   U45 : OAI21_X1 port map( B1 => n143, B2 => ENABLE, A => n175, ZN => n111);
   U46 : NAND2_X1 port map( A1 => D(20), A2 => ENABLE, ZN => n175);
   U47 : OAI21_X1 port map( B1 => n142, B2 => ENABLE, A => n174, ZN => n110);
   U48 : NAND2_X1 port map( A1 => D(21), A2 => ENABLE, ZN => n174);
   U49 : OAI21_X1 port map( B1 => n141, B2 => ENABLE, A => n173, ZN => n109);
   U50 : NAND2_X1 port map( A1 => D(22), A2 => ENABLE, ZN => n173);
   U51 : OAI21_X1 port map( B1 => n140, B2 => ENABLE, A => n172, ZN => n108);
   U52 : NAND2_X1 port map( A1 => D(23), A2 => ENABLE, ZN => n172);
   U53 : OAI21_X1 port map( B1 => n139, B2 => ENABLE, A => n171, ZN => n107);
   U54 : NAND2_X1 port map( A1 => D(24), A2 => ENABLE, ZN => n171);
   U55 : OAI21_X1 port map( B1 => n138, B2 => ENABLE, A => n170, ZN => n106);
   U56 : NAND2_X1 port map( A1 => D(25), A2 => ENABLE, ZN => n170);
   U57 : OAI21_X1 port map( B1 => n137, B2 => ENABLE, A => n169, ZN => n105);
   U58 : NAND2_X1 port map( A1 => D(26), A2 => ENABLE, ZN => n169);
   U59 : OAI21_X1 port map( B1 => n136, B2 => ENABLE, A => n168, ZN => n104);
   U60 : NAND2_X1 port map( A1 => D(27), A2 => ENABLE, ZN => n168);
   U61 : OAI21_X1 port map( B1 => n135, B2 => ENABLE, A => n167, ZN => n103);
   U62 : NAND2_X1 port map( A1 => D(28), A2 => ENABLE, ZN => n167);
   U63 : OAI21_X1 port map( B1 => n134, B2 => ENABLE, A => n166, ZN => n102);
   U64 : NAND2_X1 port map( A1 => D(29), A2 => ENABLE, ZN => n166);
   U65 : OAI21_X1 port map( B1 => n133, B2 => ENABLE, A => n165, ZN => n101);
   U66 : NAND2_X1 port map( A1 => D(30), A2 => ENABLE, ZN => n165);
   U67 : OAI21_X1 port map( B1 => n132, B2 => ENABLE, A => n164, ZN => n100);
   U68 : NAND2_X1 port map( A1 => D(31), A2 => ENABLE, ZN => n164);

end SYN_ASYNCHBEHAV;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity regFFD_NBIT32_6 is

   port( CK, RESET, ENABLE : in std_logic;  D : in std_logic_vector (31 downto 
         0);  Q : out std_logic_vector (31 downto 0));

end regFFD_NBIT32_6;

architecture SYN_ASYNCHBEHAV of regFFD_NBIT32_6 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, 
      n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, 
      n121, n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, 
      n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, 
      n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, 
      n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, 
      n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, 
      n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, 
      n193, n194, n195 : std_logic;

begin
   
   Q_reg_31_inst : DFFR_X1 port map( D => n100, CK => CK, RN => n99, Q => Q(31)
                           , QN => n132);
   Q_reg_30_inst : DFFR_X1 port map( D => n101, CK => CK, RN => n99, Q => Q(30)
                           , QN => n133);
   Q_reg_29_inst : DFFR_X1 port map( D => n102, CK => CK, RN => n99, Q => Q(29)
                           , QN => n134);
   Q_reg_28_inst : DFFR_X1 port map( D => n103, CK => CK, RN => n99, Q => Q(28)
                           , QN => n135);
   Q_reg_27_inst : DFFR_X1 port map( D => n104, CK => CK, RN => n99, Q => Q(27)
                           , QN => n136);
   Q_reg_26_inst : DFFR_X1 port map( D => n105, CK => CK, RN => n99, Q => Q(26)
                           , QN => n137);
   Q_reg_25_inst : DFFR_X1 port map( D => n106, CK => CK, RN => n99, Q => Q(25)
                           , QN => n138);
   Q_reg_24_inst : DFFR_X1 port map( D => n107, CK => CK, RN => n99, Q => Q(24)
                           , QN => n139);
   Q_reg_23_inst : DFFR_X1 port map( D => n108, CK => CK, RN => n98, Q => Q(23)
                           , QN => n140);
   Q_reg_22_inst : DFFR_X1 port map( D => n109, CK => CK, RN => n98, Q => Q(22)
                           , QN => n141);
   Q_reg_21_inst : DFFR_X1 port map( D => n110, CK => CK, RN => n98, Q => Q(21)
                           , QN => n142);
   Q_reg_20_inst : DFFR_X1 port map( D => n111, CK => CK, RN => n98, Q => Q(20)
                           , QN => n143);
   Q_reg_19_inst : DFFR_X1 port map( D => n112, CK => CK, RN => n98, Q => Q(19)
                           , QN => n144);
   Q_reg_18_inst : DFFR_X1 port map( D => n113, CK => CK, RN => n98, Q => Q(18)
                           , QN => n145);
   Q_reg_17_inst : DFFR_X1 port map( D => n114, CK => CK, RN => n98, Q => Q(17)
                           , QN => n146);
   Q_reg_16_inst : DFFR_X1 port map( D => n115, CK => CK, RN => n98, Q => Q(16)
                           , QN => n147);
   Q_reg_15_inst : DFFR_X1 port map( D => n116, CK => CK, RN => n98, Q => Q(15)
                           , QN => n148);
   Q_reg_14_inst : DFFR_X1 port map( D => n117, CK => CK, RN => n98, Q => Q(14)
                           , QN => n149);
   Q_reg_13_inst : DFFR_X1 port map( D => n118, CK => CK, RN => n98, Q => Q(13)
                           , QN => n150);
   Q_reg_12_inst : DFFR_X1 port map( D => n119, CK => CK, RN => n98, Q => Q(12)
                           , QN => n151);
   Q_reg_11_inst : DFFR_X1 port map( D => n120, CK => CK, RN => n97, Q => Q(11)
                           , QN => n152);
   Q_reg_10_inst : DFFR_X1 port map( D => n121, CK => CK, RN => n97, Q => Q(10)
                           , QN => n153);
   Q_reg_9_inst : DFFR_X1 port map( D => n122, CK => CK, RN => n97, Q => Q(9), 
                           QN => n154);
   Q_reg_8_inst : DFFR_X1 port map( D => n123, CK => CK, RN => n97, Q => Q(8), 
                           QN => n155);
   Q_reg_7_inst : DFFR_X1 port map( D => n124, CK => CK, RN => n97, Q => Q(7), 
                           QN => n156);
   Q_reg_6_inst : DFFR_X1 port map( D => n125, CK => CK, RN => n97, Q => Q(6), 
                           QN => n157);
   Q_reg_5_inst : DFFR_X1 port map( D => n126, CK => CK, RN => n97, Q => Q(5), 
                           QN => n158);
   Q_reg_4_inst : DFFR_X1 port map( D => n127, CK => CK, RN => n97, Q => Q(4), 
                           QN => n159);
   Q_reg_3_inst : DFFR_X1 port map( D => n128, CK => CK, RN => n97, Q => Q(3), 
                           QN => n160);
   Q_reg_2_inst : DFFR_X1 port map( D => n129, CK => CK, RN => n97, Q => Q(2), 
                           QN => n161);
   Q_reg_1_inst : DFFR_X1 port map( D => n130, CK => CK, RN => n97, Q => Q(1), 
                           QN => n162);
   Q_reg_0_inst : DFFR_X1 port map( D => n131, CK => CK, RN => n97, Q => Q(0), 
                           QN => n163);
   U2 : BUF_X1 port map( A => RESET, Z => n97);
   U3 : BUF_X1 port map( A => RESET, Z => n98);
   U4 : BUF_X1 port map( A => RESET, Z => n99);
   U5 : OAI21_X1 port map( B1 => n147, B2 => ENABLE, A => n179, ZN => n115);
   U6 : NAND2_X1 port map( A1 => D(16), A2 => ENABLE, ZN => n179);
   U7 : OAI21_X1 port map( B1 => n146, B2 => ENABLE, A => n178, ZN => n114);
   U8 : NAND2_X1 port map( A1 => D(17), A2 => ENABLE, ZN => n178);
   U9 : OAI21_X1 port map( B1 => n145, B2 => ENABLE, A => n177, ZN => n113);
   U10 : NAND2_X1 port map( A1 => D(18), A2 => ENABLE, ZN => n177);
   U11 : OAI21_X1 port map( B1 => n144, B2 => ENABLE, A => n176, ZN => n112);
   U12 : NAND2_X1 port map( A1 => D(19), A2 => ENABLE, ZN => n176);
   U13 : OAI21_X1 port map( B1 => n143, B2 => ENABLE, A => n175, ZN => n111);
   U14 : NAND2_X1 port map( A1 => D(20), A2 => ENABLE, ZN => n175);
   U15 : OAI21_X1 port map( B1 => n142, B2 => ENABLE, A => n174, ZN => n110);
   U16 : NAND2_X1 port map( A1 => D(21), A2 => ENABLE, ZN => n174);
   U17 : OAI21_X1 port map( B1 => n141, B2 => ENABLE, A => n173, ZN => n109);
   U18 : NAND2_X1 port map( A1 => D(22), A2 => ENABLE, ZN => n173);
   U19 : OAI21_X1 port map( B1 => n140, B2 => ENABLE, A => n172, ZN => n108);
   U20 : NAND2_X1 port map( A1 => D(23), A2 => ENABLE, ZN => n172);
   U21 : OAI21_X1 port map( B1 => n139, B2 => ENABLE, A => n171, ZN => n107);
   U22 : NAND2_X1 port map( A1 => D(24), A2 => ENABLE, ZN => n171);
   U23 : OAI21_X1 port map( B1 => n138, B2 => ENABLE, A => n170, ZN => n106);
   U24 : NAND2_X1 port map( A1 => D(25), A2 => ENABLE, ZN => n170);
   U25 : OAI21_X1 port map( B1 => n137, B2 => ENABLE, A => n169, ZN => n105);
   U26 : NAND2_X1 port map( A1 => D(26), A2 => ENABLE, ZN => n169);
   U27 : OAI21_X1 port map( B1 => n136, B2 => ENABLE, A => n168, ZN => n104);
   U28 : NAND2_X1 port map( A1 => D(27), A2 => ENABLE, ZN => n168);
   U29 : OAI21_X1 port map( B1 => n135, B2 => ENABLE, A => n167, ZN => n103);
   U30 : NAND2_X1 port map( A1 => D(28), A2 => ENABLE, ZN => n167);
   U31 : OAI21_X1 port map( B1 => n134, B2 => ENABLE, A => n166, ZN => n102);
   U32 : NAND2_X1 port map( A1 => D(29), A2 => ENABLE, ZN => n166);
   U33 : OAI21_X1 port map( B1 => n133, B2 => ENABLE, A => n165, ZN => n101);
   U34 : NAND2_X1 port map( A1 => D(30), A2 => ENABLE, ZN => n165);
   U35 : OAI21_X1 port map( B1 => n132, B2 => ENABLE, A => n164, ZN => n100);
   U36 : NAND2_X1 port map( A1 => D(31), A2 => ENABLE, ZN => n164);
   U37 : OAI21_X1 port map( B1 => n163, B2 => ENABLE, A => n195, ZN => n131);
   U38 : NAND2_X1 port map( A1 => ENABLE, A2 => D(0), ZN => n195);
   U39 : OAI21_X1 port map( B1 => n162, B2 => ENABLE, A => n194, ZN => n130);
   U40 : NAND2_X1 port map( A1 => D(1), A2 => ENABLE, ZN => n194);
   U41 : OAI21_X1 port map( B1 => n161, B2 => ENABLE, A => n193, ZN => n129);
   U42 : NAND2_X1 port map( A1 => D(2), A2 => ENABLE, ZN => n193);
   U43 : OAI21_X1 port map( B1 => n160, B2 => ENABLE, A => n192, ZN => n128);
   U44 : NAND2_X1 port map( A1 => D(3), A2 => ENABLE, ZN => n192);
   U45 : OAI21_X1 port map( B1 => n159, B2 => ENABLE, A => n191, ZN => n127);
   U46 : NAND2_X1 port map( A1 => D(4), A2 => ENABLE, ZN => n191);
   U47 : OAI21_X1 port map( B1 => n158, B2 => ENABLE, A => n190, ZN => n126);
   U48 : NAND2_X1 port map( A1 => D(5), A2 => ENABLE, ZN => n190);
   U49 : OAI21_X1 port map( B1 => n157, B2 => ENABLE, A => n189, ZN => n125);
   U50 : NAND2_X1 port map( A1 => D(6), A2 => ENABLE, ZN => n189);
   U51 : OAI21_X1 port map( B1 => n156, B2 => ENABLE, A => n188, ZN => n124);
   U52 : NAND2_X1 port map( A1 => D(7), A2 => ENABLE, ZN => n188);
   U53 : OAI21_X1 port map( B1 => n155, B2 => ENABLE, A => n187, ZN => n123);
   U54 : NAND2_X1 port map( A1 => D(8), A2 => ENABLE, ZN => n187);
   U55 : OAI21_X1 port map( B1 => n154, B2 => ENABLE, A => n186, ZN => n122);
   U56 : NAND2_X1 port map( A1 => D(9), A2 => ENABLE, ZN => n186);
   U57 : OAI21_X1 port map( B1 => n153, B2 => ENABLE, A => n185, ZN => n121);
   U58 : NAND2_X1 port map( A1 => D(10), A2 => ENABLE, ZN => n185);
   U59 : OAI21_X1 port map( B1 => n152, B2 => ENABLE, A => n184, ZN => n120);
   U60 : NAND2_X1 port map( A1 => D(11), A2 => ENABLE, ZN => n184);
   U61 : OAI21_X1 port map( B1 => n151, B2 => ENABLE, A => n183, ZN => n119);
   U62 : NAND2_X1 port map( A1 => D(12), A2 => ENABLE, ZN => n183);
   U63 : OAI21_X1 port map( B1 => n150, B2 => ENABLE, A => n182, ZN => n118);
   U64 : NAND2_X1 port map( A1 => D(13), A2 => ENABLE, ZN => n182);
   U65 : OAI21_X1 port map( B1 => n149, B2 => ENABLE, A => n181, ZN => n117);
   U66 : NAND2_X1 port map( A1 => D(14), A2 => ENABLE, ZN => n181);
   U67 : OAI21_X1 port map( B1 => n148, B2 => ENABLE, A => n180, ZN => n116);
   U68 : NAND2_X1 port map( A1 => D(15), A2 => ENABLE, ZN => n180);

end SYN_ASYNCHBEHAV;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity regFFD_NBIT32_5 is

   port( CK, RESET, ENABLE : in std_logic;  D : in std_logic_vector (31 downto 
         0);  Q : out std_logic_vector (31 downto 0));

end regFFD_NBIT32_5;

architecture SYN_ASYNCHBEHAV of regFFD_NBIT32_5 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, 
      n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, 
      n121, n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, 
      n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, 
      n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, 
      n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, 
      n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, 
      n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, 
      n193, n194, n195 : std_logic;

begin
   
   Q_reg_31_inst : DFFR_X1 port map( D => n100, CK => CK, RN => n99, Q => Q(31)
                           , QN => n132);
   Q_reg_30_inst : DFFR_X1 port map( D => n101, CK => CK, RN => n99, Q => Q(30)
                           , QN => n133);
   Q_reg_29_inst : DFFR_X1 port map( D => n102, CK => CK, RN => n99, Q => Q(29)
                           , QN => n134);
   Q_reg_28_inst : DFFR_X1 port map( D => n103, CK => CK, RN => n99, Q => Q(28)
                           , QN => n135);
   Q_reg_27_inst : DFFR_X1 port map( D => n104, CK => CK, RN => n99, Q => Q(27)
                           , QN => n136);
   Q_reg_26_inst : DFFR_X1 port map( D => n105, CK => CK, RN => n99, Q => Q(26)
                           , QN => n137);
   Q_reg_25_inst : DFFR_X1 port map( D => n106, CK => CK, RN => n99, Q => Q(25)
                           , QN => n138);
   Q_reg_24_inst : DFFR_X1 port map( D => n107, CK => CK, RN => n99, Q => Q(24)
                           , QN => n139);
   Q_reg_23_inst : DFFR_X1 port map( D => n108, CK => CK, RN => n98, Q => Q(23)
                           , QN => n140);
   Q_reg_22_inst : DFFR_X1 port map( D => n109, CK => CK, RN => n98, Q => Q(22)
                           , QN => n141);
   Q_reg_21_inst : DFFR_X1 port map( D => n110, CK => CK, RN => n98, Q => Q(21)
                           , QN => n142);
   Q_reg_20_inst : DFFR_X1 port map( D => n111, CK => CK, RN => n98, Q => Q(20)
                           , QN => n143);
   Q_reg_19_inst : DFFR_X1 port map( D => n112, CK => CK, RN => n98, Q => Q(19)
                           , QN => n144);
   Q_reg_18_inst : DFFR_X1 port map( D => n113, CK => CK, RN => n98, Q => Q(18)
                           , QN => n145);
   Q_reg_17_inst : DFFR_X1 port map( D => n114, CK => CK, RN => n98, Q => Q(17)
                           , QN => n146);
   Q_reg_16_inst : DFFR_X1 port map( D => n115, CK => CK, RN => n98, Q => Q(16)
                           , QN => n147);
   Q_reg_15_inst : DFFR_X1 port map( D => n116, CK => CK, RN => n98, Q => Q(15)
                           , QN => n148);
   Q_reg_14_inst : DFFR_X1 port map( D => n117, CK => CK, RN => n98, Q => Q(14)
                           , QN => n149);
   Q_reg_13_inst : DFFR_X1 port map( D => n118, CK => CK, RN => n98, Q => Q(13)
                           , QN => n150);
   Q_reg_12_inst : DFFR_X1 port map( D => n119, CK => CK, RN => n98, Q => Q(12)
                           , QN => n151);
   Q_reg_11_inst : DFFR_X1 port map( D => n120, CK => CK, RN => n97, Q => Q(11)
                           , QN => n152);
   Q_reg_10_inst : DFFR_X1 port map( D => n121, CK => CK, RN => n97, Q => Q(10)
                           , QN => n153);
   Q_reg_9_inst : DFFR_X1 port map( D => n122, CK => CK, RN => n97, Q => Q(9), 
                           QN => n154);
   Q_reg_8_inst : DFFR_X1 port map( D => n123, CK => CK, RN => n97, Q => Q(8), 
                           QN => n155);
   Q_reg_7_inst : DFFR_X1 port map( D => n124, CK => CK, RN => n97, Q => Q(7), 
                           QN => n156);
   Q_reg_6_inst : DFFR_X1 port map( D => n125, CK => CK, RN => n97, Q => Q(6), 
                           QN => n157);
   Q_reg_5_inst : DFFR_X1 port map( D => n126, CK => CK, RN => n97, Q => Q(5), 
                           QN => n158);
   Q_reg_4_inst : DFFR_X1 port map( D => n127, CK => CK, RN => n97, Q => Q(4), 
                           QN => n159);
   Q_reg_3_inst : DFFR_X1 port map( D => n128, CK => CK, RN => n97, Q => Q(3), 
                           QN => n160);
   Q_reg_2_inst : DFFR_X1 port map( D => n129, CK => CK, RN => n97, Q => Q(2), 
                           QN => n161);
   Q_reg_1_inst : DFFR_X1 port map( D => n130, CK => CK, RN => n97, Q => Q(1), 
                           QN => n162);
   Q_reg_0_inst : DFFR_X1 port map( D => n131, CK => CK, RN => n97, Q => Q(0), 
                           QN => n163);
   U2 : BUF_X1 port map( A => RESET, Z => n97);
   U3 : BUF_X1 port map( A => RESET, Z => n98);
   U4 : BUF_X1 port map( A => RESET, Z => n99);
   U5 : OAI21_X1 port map( B1 => n163, B2 => ENABLE, A => n195, ZN => n131);
   U6 : NAND2_X1 port map( A1 => ENABLE, A2 => D(0), ZN => n195);
   U7 : OAI21_X1 port map( B1 => n162, B2 => ENABLE, A => n194, ZN => n130);
   U8 : NAND2_X1 port map( A1 => D(1), A2 => ENABLE, ZN => n194);
   U9 : OAI21_X1 port map( B1 => n161, B2 => ENABLE, A => n193, ZN => n129);
   U10 : NAND2_X1 port map( A1 => D(2), A2 => ENABLE, ZN => n193);
   U11 : OAI21_X1 port map( B1 => n160, B2 => ENABLE, A => n192, ZN => n128);
   U12 : NAND2_X1 port map( A1 => D(3), A2 => ENABLE, ZN => n192);
   U13 : OAI21_X1 port map( B1 => n159, B2 => ENABLE, A => n191, ZN => n127);
   U14 : NAND2_X1 port map( A1 => D(4), A2 => ENABLE, ZN => n191);
   U15 : OAI21_X1 port map( B1 => n158, B2 => ENABLE, A => n190, ZN => n126);
   U16 : NAND2_X1 port map( A1 => D(5), A2 => ENABLE, ZN => n190);
   U17 : OAI21_X1 port map( B1 => n157, B2 => ENABLE, A => n189, ZN => n125);
   U18 : NAND2_X1 port map( A1 => D(6), A2 => ENABLE, ZN => n189);
   U19 : OAI21_X1 port map( B1 => n156, B2 => ENABLE, A => n188, ZN => n124);
   U20 : NAND2_X1 port map( A1 => D(7), A2 => ENABLE, ZN => n188);
   U21 : OAI21_X1 port map( B1 => n155, B2 => ENABLE, A => n187, ZN => n123);
   U22 : NAND2_X1 port map( A1 => D(8), A2 => ENABLE, ZN => n187);
   U23 : OAI21_X1 port map( B1 => n154, B2 => ENABLE, A => n186, ZN => n122);
   U24 : NAND2_X1 port map( A1 => D(9), A2 => ENABLE, ZN => n186);
   U25 : OAI21_X1 port map( B1 => n153, B2 => ENABLE, A => n185, ZN => n121);
   U26 : NAND2_X1 port map( A1 => D(10), A2 => ENABLE, ZN => n185);
   U27 : OAI21_X1 port map( B1 => n152, B2 => ENABLE, A => n184, ZN => n120);
   U28 : NAND2_X1 port map( A1 => D(11), A2 => ENABLE, ZN => n184);
   U29 : OAI21_X1 port map( B1 => n151, B2 => ENABLE, A => n183, ZN => n119);
   U30 : NAND2_X1 port map( A1 => D(12), A2 => ENABLE, ZN => n183);
   U31 : OAI21_X1 port map( B1 => n150, B2 => ENABLE, A => n182, ZN => n118);
   U32 : NAND2_X1 port map( A1 => D(13), A2 => ENABLE, ZN => n182);
   U33 : OAI21_X1 port map( B1 => n149, B2 => ENABLE, A => n181, ZN => n117);
   U34 : NAND2_X1 port map( A1 => D(14), A2 => ENABLE, ZN => n181);
   U35 : OAI21_X1 port map( B1 => n148, B2 => ENABLE, A => n180, ZN => n116);
   U36 : NAND2_X1 port map( A1 => D(15), A2 => ENABLE, ZN => n180);
   U37 : OAI21_X1 port map( B1 => n147, B2 => ENABLE, A => n179, ZN => n115);
   U38 : NAND2_X1 port map( A1 => D(16), A2 => ENABLE, ZN => n179);
   U39 : OAI21_X1 port map( B1 => n146, B2 => ENABLE, A => n178, ZN => n114);
   U40 : NAND2_X1 port map( A1 => D(17), A2 => ENABLE, ZN => n178);
   U41 : OAI21_X1 port map( B1 => n145, B2 => ENABLE, A => n177, ZN => n113);
   U42 : NAND2_X1 port map( A1 => D(18), A2 => ENABLE, ZN => n177);
   U43 : OAI21_X1 port map( B1 => n144, B2 => ENABLE, A => n176, ZN => n112);
   U44 : NAND2_X1 port map( A1 => D(19), A2 => ENABLE, ZN => n176);
   U45 : OAI21_X1 port map( B1 => n143, B2 => ENABLE, A => n175, ZN => n111);
   U46 : NAND2_X1 port map( A1 => D(20), A2 => ENABLE, ZN => n175);
   U47 : OAI21_X1 port map( B1 => n142, B2 => ENABLE, A => n174, ZN => n110);
   U48 : NAND2_X1 port map( A1 => D(21), A2 => ENABLE, ZN => n174);
   U49 : OAI21_X1 port map( B1 => n141, B2 => ENABLE, A => n173, ZN => n109);
   U50 : NAND2_X1 port map( A1 => D(22), A2 => ENABLE, ZN => n173);
   U51 : OAI21_X1 port map( B1 => n140, B2 => ENABLE, A => n172, ZN => n108);
   U52 : NAND2_X1 port map( A1 => D(23), A2 => ENABLE, ZN => n172);
   U53 : OAI21_X1 port map( B1 => n139, B2 => ENABLE, A => n171, ZN => n107);
   U54 : NAND2_X1 port map( A1 => D(24), A2 => ENABLE, ZN => n171);
   U55 : OAI21_X1 port map( B1 => n138, B2 => ENABLE, A => n170, ZN => n106);
   U56 : NAND2_X1 port map( A1 => D(25), A2 => ENABLE, ZN => n170);
   U57 : OAI21_X1 port map( B1 => n137, B2 => ENABLE, A => n169, ZN => n105);
   U58 : NAND2_X1 port map( A1 => D(26), A2 => ENABLE, ZN => n169);
   U59 : OAI21_X1 port map( B1 => n136, B2 => ENABLE, A => n168, ZN => n104);
   U60 : NAND2_X1 port map( A1 => D(27), A2 => ENABLE, ZN => n168);
   U61 : OAI21_X1 port map( B1 => n135, B2 => ENABLE, A => n167, ZN => n103);
   U62 : NAND2_X1 port map( A1 => D(28), A2 => ENABLE, ZN => n167);
   U63 : OAI21_X1 port map( B1 => n134, B2 => ENABLE, A => n166, ZN => n102);
   U64 : NAND2_X1 port map( A1 => D(29), A2 => ENABLE, ZN => n166);
   U65 : OAI21_X1 port map( B1 => n133, B2 => ENABLE, A => n165, ZN => n101);
   U66 : NAND2_X1 port map( A1 => D(30), A2 => ENABLE, ZN => n165);
   U67 : OAI21_X1 port map( B1 => n132, B2 => ENABLE, A => n164, ZN => n100);
   U68 : NAND2_X1 port map( A1 => D(31), A2 => ENABLE, ZN => n164);

end SYN_ASYNCHBEHAV;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity regFFD_NBIT32_4 is

   port( CK, RESET, ENABLE : in std_logic;  D : in std_logic_vector (31 downto 
         0);  Q : out std_logic_vector (31 downto 0));

end regFFD_NBIT32_4;

architecture SYN_ASYNCHBEHAV of regFFD_NBIT32_4 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, 
      n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, 
      n121, n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, 
      n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, 
      n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, 
      n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, 
      n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, 
      n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, 
      n193, n194, n195 : std_logic;

begin
   
   Q_reg_31_inst : DFFR_X1 port map( D => n100, CK => CK, RN => n99, Q => Q(31)
                           , QN => n132);
   Q_reg_30_inst : DFFR_X1 port map( D => n101, CK => CK, RN => n99, Q => Q(30)
                           , QN => n133);
   Q_reg_29_inst : DFFR_X1 port map( D => n102, CK => CK, RN => n99, Q => Q(29)
                           , QN => n134);
   Q_reg_28_inst : DFFR_X1 port map( D => n103, CK => CK, RN => n99, Q => Q(28)
                           , QN => n135);
   Q_reg_27_inst : DFFR_X1 port map( D => n104, CK => CK, RN => n99, Q => Q(27)
                           , QN => n136);
   Q_reg_26_inst : DFFR_X1 port map( D => n105, CK => CK, RN => n99, Q => Q(26)
                           , QN => n137);
   Q_reg_25_inst : DFFR_X1 port map( D => n106, CK => CK, RN => n99, Q => Q(25)
                           , QN => n138);
   Q_reg_24_inst : DFFR_X1 port map( D => n107, CK => CK, RN => n99, Q => Q(24)
                           , QN => n139);
   Q_reg_23_inst : DFFR_X1 port map( D => n108, CK => CK, RN => n98, Q => Q(23)
                           , QN => n140);
   Q_reg_22_inst : DFFR_X1 port map( D => n109, CK => CK, RN => n98, Q => Q(22)
                           , QN => n141);
   Q_reg_21_inst : DFFR_X1 port map( D => n110, CK => CK, RN => n98, Q => Q(21)
                           , QN => n142);
   Q_reg_20_inst : DFFR_X1 port map( D => n111, CK => CK, RN => n98, Q => Q(20)
                           , QN => n143);
   Q_reg_19_inst : DFFR_X1 port map( D => n112, CK => CK, RN => n98, Q => Q(19)
                           , QN => n144);
   Q_reg_18_inst : DFFR_X1 port map( D => n113, CK => CK, RN => n98, Q => Q(18)
                           , QN => n145);
   Q_reg_17_inst : DFFR_X1 port map( D => n114, CK => CK, RN => n98, Q => Q(17)
                           , QN => n146);
   Q_reg_16_inst : DFFR_X1 port map( D => n115, CK => CK, RN => n98, Q => Q(16)
                           , QN => n147);
   Q_reg_15_inst : DFFR_X1 port map( D => n116, CK => CK, RN => n98, Q => Q(15)
                           , QN => n148);
   Q_reg_14_inst : DFFR_X1 port map( D => n117, CK => CK, RN => n98, Q => Q(14)
                           , QN => n149);
   Q_reg_13_inst : DFFR_X1 port map( D => n118, CK => CK, RN => n98, Q => Q(13)
                           , QN => n150);
   Q_reg_12_inst : DFFR_X1 port map( D => n119, CK => CK, RN => n98, Q => Q(12)
                           , QN => n151);
   Q_reg_11_inst : DFFR_X1 port map( D => n120, CK => CK, RN => n97, Q => Q(11)
                           , QN => n152);
   Q_reg_10_inst : DFFR_X1 port map( D => n121, CK => CK, RN => n97, Q => Q(10)
                           , QN => n153);
   Q_reg_9_inst : DFFR_X1 port map( D => n122, CK => CK, RN => n97, Q => Q(9), 
                           QN => n154);
   Q_reg_8_inst : DFFR_X1 port map( D => n123, CK => CK, RN => n97, Q => Q(8), 
                           QN => n155);
   Q_reg_7_inst : DFFR_X1 port map( D => n124, CK => CK, RN => n97, Q => Q(7), 
                           QN => n156);
   Q_reg_6_inst : DFFR_X1 port map( D => n125, CK => CK, RN => n97, Q => Q(6), 
                           QN => n157);
   Q_reg_5_inst : DFFR_X1 port map( D => n126, CK => CK, RN => n97, Q => Q(5), 
                           QN => n158);
   Q_reg_4_inst : DFFR_X1 port map( D => n127, CK => CK, RN => n97, Q => Q(4), 
                           QN => n159);
   Q_reg_3_inst : DFFR_X1 port map( D => n128, CK => CK, RN => n97, Q => Q(3), 
                           QN => n160);
   Q_reg_2_inst : DFFR_X1 port map( D => n129, CK => CK, RN => n97, Q => Q(2), 
                           QN => n161);
   Q_reg_1_inst : DFFR_X1 port map( D => n130, CK => CK, RN => n97, Q => Q(1), 
                           QN => n162);
   Q_reg_0_inst : DFFR_X1 port map( D => n131, CK => CK, RN => n97, Q => Q(0), 
                           QN => n163);
   U2 : BUF_X1 port map( A => RESET, Z => n97);
   U3 : BUF_X1 port map( A => RESET, Z => n98);
   U4 : BUF_X1 port map( A => RESET, Z => n99);
   U5 : OAI21_X1 port map( B1 => n163, B2 => ENABLE, A => n195, ZN => n131);
   U6 : NAND2_X1 port map( A1 => ENABLE, A2 => D(0), ZN => n195);
   U7 : OAI21_X1 port map( B1 => n162, B2 => ENABLE, A => n194, ZN => n130);
   U8 : NAND2_X1 port map( A1 => D(1), A2 => ENABLE, ZN => n194);
   U9 : OAI21_X1 port map( B1 => n161, B2 => ENABLE, A => n193, ZN => n129);
   U10 : NAND2_X1 port map( A1 => D(2), A2 => ENABLE, ZN => n193);
   U11 : OAI21_X1 port map( B1 => n160, B2 => ENABLE, A => n192, ZN => n128);
   U12 : NAND2_X1 port map( A1 => D(3), A2 => ENABLE, ZN => n192);
   U13 : OAI21_X1 port map( B1 => n159, B2 => ENABLE, A => n191, ZN => n127);
   U14 : NAND2_X1 port map( A1 => D(4), A2 => ENABLE, ZN => n191);
   U15 : OAI21_X1 port map( B1 => n158, B2 => ENABLE, A => n190, ZN => n126);
   U16 : NAND2_X1 port map( A1 => D(5), A2 => ENABLE, ZN => n190);
   U17 : OAI21_X1 port map( B1 => n157, B2 => ENABLE, A => n189, ZN => n125);
   U18 : NAND2_X1 port map( A1 => D(6), A2 => ENABLE, ZN => n189);
   U19 : OAI21_X1 port map( B1 => n156, B2 => ENABLE, A => n188, ZN => n124);
   U20 : NAND2_X1 port map( A1 => D(7), A2 => ENABLE, ZN => n188);
   U21 : OAI21_X1 port map( B1 => n155, B2 => ENABLE, A => n187, ZN => n123);
   U22 : NAND2_X1 port map( A1 => D(8), A2 => ENABLE, ZN => n187);
   U23 : OAI21_X1 port map( B1 => n154, B2 => ENABLE, A => n186, ZN => n122);
   U24 : NAND2_X1 port map( A1 => D(9), A2 => ENABLE, ZN => n186);
   U25 : OAI21_X1 port map( B1 => n153, B2 => ENABLE, A => n185, ZN => n121);
   U26 : NAND2_X1 port map( A1 => D(10), A2 => ENABLE, ZN => n185);
   U27 : OAI21_X1 port map( B1 => n152, B2 => ENABLE, A => n184, ZN => n120);
   U28 : NAND2_X1 port map( A1 => D(11), A2 => ENABLE, ZN => n184);
   U29 : OAI21_X1 port map( B1 => n151, B2 => ENABLE, A => n183, ZN => n119);
   U30 : NAND2_X1 port map( A1 => D(12), A2 => ENABLE, ZN => n183);
   U31 : OAI21_X1 port map( B1 => n150, B2 => ENABLE, A => n182, ZN => n118);
   U32 : NAND2_X1 port map( A1 => D(13), A2 => ENABLE, ZN => n182);
   U33 : OAI21_X1 port map( B1 => n149, B2 => ENABLE, A => n181, ZN => n117);
   U34 : NAND2_X1 port map( A1 => D(14), A2 => ENABLE, ZN => n181);
   U35 : OAI21_X1 port map( B1 => n148, B2 => ENABLE, A => n180, ZN => n116);
   U36 : NAND2_X1 port map( A1 => D(15), A2 => ENABLE, ZN => n180);
   U37 : OAI21_X1 port map( B1 => n147, B2 => ENABLE, A => n179, ZN => n115);
   U38 : NAND2_X1 port map( A1 => D(16), A2 => ENABLE, ZN => n179);
   U39 : OAI21_X1 port map( B1 => n146, B2 => ENABLE, A => n178, ZN => n114);
   U40 : NAND2_X1 port map( A1 => D(17), A2 => ENABLE, ZN => n178);
   U41 : OAI21_X1 port map( B1 => n145, B2 => ENABLE, A => n177, ZN => n113);
   U42 : NAND2_X1 port map( A1 => D(18), A2 => ENABLE, ZN => n177);
   U43 : OAI21_X1 port map( B1 => n144, B2 => ENABLE, A => n176, ZN => n112);
   U44 : NAND2_X1 port map( A1 => D(19), A2 => ENABLE, ZN => n176);
   U45 : OAI21_X1 port map( B1 => n143, B2 => ENABLE, A => n175, ZN => n111);
   U46 : NAND2_X1 port map( A1 => D(20), A2 => ENABLE, ZN => n175);
   U47 : OAI21_X1 port map( B1 => n142, B2 => ENABLE, A => n174, ZN => n110);
   U48 : NAND2_X1 port map( A1 => D(21), A2 => ENABLE, ZN => n174);
   U49 : OAI21_X1 port map( B1 => n141, B2 => ENABLE, A => n173, ZN => n109);
   U50 : NAND2_X1 port map( A1 => D(22), A2 => ENABLE, ZN => n173);
   U51 : OAI21_X1 port map( B1 => n140, B2 => ENABLE, A => n172, ZN => n108);
   U52 : NAND2_X1 port map( A1 => D(23), A2 => ENABLE, ZN => n172);
   U53 : OAI21_X1 port map( B1 => n139, B2 => ENABLE, A => n171, ZN => n107);
   U54 : NAND2_X1 port map( A1 => D(24), A2 => ENABLE, ZN => n171);
   U55 : OAI21_X1 port map( B1 => n138, B2 => ENABLE, A => n170, ZN => n106);
   U56 : NAND2_X1 port map( A1 => D(25), A2 => ENABLE, ZN => n170);
   U57 : OAI21_X1 port map( B1 => n137, B2 => ENABLE, A => n169, ZN => n105);
   U58 : NAND2_X1 port map( A1 => D(26), A2 => ENABLE, ZN => n169);
   U59 : OAI21_X1 port map( B1 => n136, B2 => ENABLE, A => n168, ZN => n104);
   U60 : NAND2_X1 port map( A1 => D(27), A2 => ENABLE, ZN => n168);
   U61 : OAI21_X1 port map( B1 => n135, B2 => ENABLE, A => n167, ZN => n103);
   U62 : NAND2_X1 port map( A1 => D(28), A2 => ENABLE, ZN => n167);
   U63 : OAI21_X1 port map( B1 => n134, B2 => ENABLE, A => n166, ZN => n102);
   U64 : NAND2_X1 port map( A1 => D(29), A2 => ENABLE, ZN => n166);
   U65 : OAI21_X1 port map( B1 => n133, B2 => ENABLE, A => n165, ZN => n101);
   U66 : NAND2_X1 port map( A1 => D(30), A2 => ENABLE, ZN => n165);
   U67 : OAI21_X1 port map( B1 => n132, B2 => ENABLE, A => n164, ZN => n100);
   U68 : NAND2_X1 port map( A1 => D(31), A2 => ENABLE, ZN => n164);

end SYN_ASYNCHBEHAV;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity regFFD_NBIT32_3 is

   port( CK, RESET, ENABLE : in std_logic;  D : in std_logic_vector (31 downto 
         0);  Q : out std_logic_vector (31 downto 0));

end regFFD_NBIT32_3;

architecture SYN_ASYNCHBEHAV of regFFD_NBIT32_3 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, 
      n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, 
      n121, n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, 
      n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, 
      n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, 
      n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, 
      n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, 
      n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, 
      n193, n194, n195 : std_logic;

begin
   
   Q_reg_31_inst : DFFR_X1 port map( D => n100, CK => CK, RN => n99, Q => Q(31)
                           , QN => n132);
   Q_reg_30_inst : DFFR_X1 port map( D => n101, CK => CK, RN => n99, Q => Q(30)
                           , QN => n133);
   Q_reg_29_inst : DFFR_X1 port map( D => n102, CK => CK, RN => n99, Q => Q(29)
                           , QN => n134);
   Q_reg_28_inst : DFFR_X1 port map( D => n103, CK => CK, RN => n99, Q => Q(28)
                           , QN => n135);
   Q_reg_27_inst : DFFR_X1 port map( D => n104, CK => CK, RN => n99, Q => Q(27)
                           , QN => n136);
   Q_reg_26_inst : DFFR_X1 port map( D => n105, CK => CK, RN => n99, Q => Q(26)
                           , QN => n137);
   Q_reg_25_inst : DFFR_X1 port map( D => n106, CK => CK, RN => n99, Q => Q(25)
                           , QN => n138);
   Q_reg_24_inst : DFFR_X1 port map( D => n107, CK => CK, RN => n99, Q => Q(24)
                           , QN => n139);
   Q_reg_23_inst : DFFR_X1 port map( D => n108, CK => CK, RN => n98, Q => Q(23)
                           , QN => n140);
   Q_reg_22_inst : DFFR_X1 port map( D => n109, CK => CK, RN => n98, Q => Q(22)
                           , QN => n141);
   Q_reg_21_inst : DFFR_X1 port map( D => n110, CK => CK, RN => n98, Q => Q(21)
                           , QN => n142);
   Q_reg_20_inst : DFFR_X1 port map( D => n111, CK => CK, RN => n98, Q => Q(20)
                           , QN => n143);
   Q_reg_19_inst : DFFR_X1 port map( D => n112, CK => CK, RN => n98, Q => Q(19)
                           , QN => n144);
   Q_reg_18_inst : DFFR_X1 port map( D => n113, CK => CK, RN => n98, Q => Q(18)
                           , QN => n145);
   Q_reg_17_inst : DFFR_X1 port map( D => n114, CK => CK, RN => n98, Q => Q(17)
                           , QN => n146);
   Q_reg_16_inst : DFFR_X1 port map( D => n115, CK => CK, RN => n98, Q => Q(16)
                           , QN => n147);
   Q_reg_15_inst : DFFR_X1 port map( D => n116, CK => CK, RN => n98, Q => Q(15)
                           , QN => n148);
   Q_reg_14_inst : DFFR_X1 port map( D => n117, CK => CK, RN => n98, Q => Q(14)
                           , QN => n149);
   Q_reg_13_inst : DFFR_X1 port map( D => n118, CK => CK, RN => n98, Q => Q(13)
                           , QN => n150);
   Q_reg_12_inst : DFFR_X1 port map( D => n119, CK => CK, RN => n98, Q => Q(12)
                           , QN => n151);
   Q_reg_11_inst : DFFR_X1 port map( D => n120, CK => CK, RN => n97, Q => Q(11)
                           , QN => n152);
   Q_reg_10_inst : DFFR_X1 port map( D => n121, CK => CK, RN => n97, Q => Q(10)
                           , QN => n153);
   Q_reg_9_inst : DFFR_X1 port map( D => n122, CK => CK, RN => n97, Q => Q(9), 
                           QN => n154);
   Q_reg_8_inst : DFFR_X1 port map( D => n123, CK => CK, RN => n97, Q => Q(8), 
                           QN => n155);
   Q_reg_7_inst : DFFR_X1 port map( D => n124, CK => CK, RN => n97, Q => Q(7), 
                           QN => n156);
   Q_reg_6_inst : DFFR_X1 port map( D => n125, CK => CK, RN => n97, Q => Q(6), 
                           QN => n157);
   Q_reg_5_inst : DFFR_X1 port map( D => n126, CK => CK, RN => n97, Q => Q(5), 
                           QN => n158);
   Q_reg_4_inst : DFFR_X1 port map( D => n127, CK => CK, RN => n97, Q => Q(4), 
                           QN => n159);
   Q_reg_3_inst : DFFR_X1 port map( D => n128, CK => CK, RN => n97, Q => Q(3), 
                           QN => n160);
   Q_reg_2_inst : DFFR_X1 port map( D => n129, CK => CK, RN => n97, Q => Q(2), 
                           QN => n161);
   Q_reg_1_inst : DFFR_X1 port map( D => n130, CK => CK, RN => n97, Q => Q(1), 
                           QN => n162);
   Q_reg_0_inst : DFFR_X1 port map( D => n131, CK => CK, RN => n97, Q => Q(0), 
                           QN => n163);
   U2 : BUF_X1 port map( A => RESET, Z => n97);
   U3 : BUF_X1 port map( A => RESET, Z => n98);
   U4 : BUF_X1 port map( A => RESET, Z => n99);
   U5 : OAI21_X1 port map( B1 => n163, B2 => ENABLE, A => n195, ZN => n131);
   U6 : NAND2_X1 port map( A1 => ENABLE, A2 => D(0), ZN => n195);
   U7 : OAI21_X1 port map( B1 => n162, B2 => ENABLE, A => n194, ZN => n130);
   U8 : NAND2_X1 port map( A1 => D(1), A2 => ENABLE, ZN => n194);
   U9 : OAI21_X1 port map( B1 => n161, B2 => ENABLE, A => n193, ZN => n129);
   U10 : NAND2_X1 port map( A1 => D(2), A2 => ENABLE, ZN => n193);
   U11 : OAI21_X1 port map( B1 => n160, B2 => ENABLE, A => n192, ZN => n128);
   U12 : NAND2_X1 port map( A1 => D(3), A2 => ENABLE, ZN => n192);
   U13 : OAI21_X1 port map( B1 => n159, B2 => ENABLE, A => n191, ZN => n127);
   U14 : NAND2_X1 port map( A1 => D(4), A2 => ENABLE, ZN => n191);
   U15 : OAI21_X1 port map( B1 => n158, B2 => ENABLE, A => n190, ZN => n126);
   U16 : NAND2_X1 port map( A1 => D(5), A2 => ENABLE, ZN => n190);
   U17 : OAI21_X1 port map( B1 => n157, B2 => ENABLE, A => n189, ZN => n125);
   U18 : NAND2_X1 port map( A1 => D(6), A2 => ENABLE, ZN => n189);
   U19 : OAI21_X1 port map( B1 => n156, B2 => ENABLE, A => n188, ZN => n124);
   U20 : NAND2_X1 port map( A1 => D(7), A2 => ENABLE, ZN => n188);
   U21 : OAI21_X1 port map( B1 => n155, B2 => ENABLE, A => n187, ZN => n123);
   U22 : NAND2_X1 port map( A1 => D(8), A2 => ENABLE, ZN => n187);
   U23 : OAI21_X1 port map( B1 => n154, B2 => ENABLE, A => n186, ZN => n122);
   U24 : NAND2_X1 port map( A1 => D(9), A2 => ENABLE, ZN => n186);
   U25 : OAI21_X1 port map( B1 => n153, B2 => ENABLE, A => n185, ZN => n121);
   U26 : NAND2_X1 port map( A1 => D(10), A2 => ENABLE, ZN => n185);
   U27 : OAI21_X1 port map( B1 => n152, B2 => ENABLE, A => n184, ZN => n120);
   U28 : NAND2_X1 port map( A1 => D(11), A2 => ENABLE, ZN => n184);
   U29 : OAI21_X1 port map( B1 => n151, B2 => ENABLE, A => n183, ZN => n119);
   U30 : NAND2_X1 port map( A1 => D(12), A2 => ENABLE, ZN => n183);
   U31 : OAI21_X1 port map( B1 => n150, B2 => ENABLE, A => n182, ZN => n118);
   U32 : NAND2_X1 port map( A1 => D(13), A2 => ENABLE, ZN => n182);
   U33 : OAI21_X1 port map( B1 => n149, B2 => ENABLE, A => n181, ZN => n117);
   U34 : NAND2_X1 port map( A1 => D(14), A2 => ENABLE, ZN => n181);
   U35 : OAI21_X1 port map( B1 => n148, B2 => ENABLE, A => n180, ZN => n116);
   U36 : NAND2_X1 port map( A1 => D(15), A2 => ENABLE, ZN => n180);
   U37 : OAI21_X1 port map( B1 => n147, B2 => ENABLE, A => n179, ZN => n115);
   U38 : NAND2_X1 port map( A1 => D(16), A2 => ENABLE, ZN => n179);
   U39 : OAI21_X1 port map( B1 => n146, B2 => ENABLE, A => n178, ZN => n114);
   U40 : NAND2_X1 port map( A1 => D(17), A2 => ENABLE, ZN => n178);
   U41 : OAI21_X1 port map( B1 => n145, B2 => ENABLE, A => n177, ZN => n113);
   U42 : NAND2_X1 port map( A1 => D(18), A2 => ENABLE, ZN => n177);
   U43 : OAI21_X1 port map( B1 => n144, B2 => ENABLE, A => n176, ZN => n112);
   U44 : NAND2_X1 port map( A1 => D(19), A2 => ENABLE, ZN => n176);
   U45 : OAI21_X1 port map( B1 => n143, B2 => ENABLE, A => n175, ZN => n111);
   U46 : NAND2_X1 port map( A1 => D(20), A2 => ENABLE, ZN => n175);
   U47 : OAI21_X1 port map( B1 => n142, B2 => ENABLE, A => n174, ZN => n110);
   U48 : NAND2_X1 port map( A1 => D(21), A2 => ENABLE, ZN => n174);
   U49 : OAI21_X1 port map( B1 => n141, B2 => ENABLE, A => n173, ZN => n109);
   U50 : NAND2_X1 port map( A1 => D(22), A2 => ENABLE, ZN => n173);
   U51 : OAI21_X1 port map( B1 => n140, B2 => ENABLE, A => n172, ZN => n108);
   U52 : NAND2_X1 port map( A1 => D(23), A2 => ENABLE, ZN => n172);
   U53 : OAI21_X1 port map( B1 => n139, B2 => ENABLE, A => n171, ZN => n107);
   U54 : NAND2_X1 port map( A1 => D(24), A2 => ENABLE, ZN => n171);
   U55 : OAI21_X1 port map( B1 => n138, B2 => ENABLE, A => n170, ZN => n106);
   U56 : NAND2_X1 port map( A1 => D(25), A2 => ENABLE, ZN => n170);
   U57 : OAI21_X1 port map( B1 => n137, B2 => ENABLE, A => n169, ZN => n105);
   U58 : NAND2_X1 port map( A1 => D(26), A2 => ENABLE, ZN => n169);
   U59 : OAI21_X1 port map( B1 => n136, B2 => ENABLE, A => n168, ZN => n104);
   U60 : NAND2_X1 port map( A1 => D(27), A2 => ENABLE, ZN => n168);
   U61 : OAI21_X1 port map( B1 => n135, B2 => ENABLE, A => n167, ZN => n103);
   U62 : NAND2_X1 port map( A1 => D(28), A2 => ENABLE, ZN => n167);
   U63 : OAI21_X1 port map( B1 => n134, B2 => ENABLE, A => n166, ZN => n102);
   U64 : NAND2_X1 port map( A1 => D(29), A2 => ENABLE, ZN => n166);
   U65 : OAI21_X1 port map( B1 => n133, B2 => ENABLE, A => n165, ZN => n101);
   U66 : NAND2_X1 port map( A1 => D(30), A2 => ENABLE, ZN => n165);
   U67 : OAI21_X1 port map( B1 => n132, B2 => ENABLE, A => n164, ZN => n100);
   U68 : NAND2_X1 port map( A1 => D(31), A2 => ENABLE, ZN => n164);

end SYN_ASYNCHBEHAV;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity regFFD_NBIT32_2 is

   port( CK, RESET, ENABLE : in std_logic;  D : in std_logic_vector (31 downto 
         0);  Q : out std_logic_vector (31 downto 0));

end regFFD_NBIT32_2;

architecture SYN_ASYNCHBEHAV of regFFD_NBIT32_2 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, 
      n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, 
      n121, n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, 
      n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, 
      n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, 
      n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, 
      n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, 
      n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, 
      n193, n194, n195 : std_logic;

begin
   
   Q_reg_31_inst : DFFR_X1 port map( D => n100, CK => CK, RN => n99, Q => Q(31)
                           , QN => n132);
   Q_reg_30_inst : DFFR_X1 port map( D => n101, CK => CK, RN => n99, Q => Q(30)
                           , QN => n133);
   Q_reg_29_inst : DFFR_X1 port map( D => n102, CK => CK, RN => n99, Q => Q(29)
                           , QN => n134);
   Q_reg_28_inst : DFFR_X1 port map( D => n103, CK => CK, RN => n99, Q => Q(28)
                           , QN => n135);
   Q_reg_27_inst : DFFR_X1 port map( D => n104, CK => CK, RN => n99, Q => Q(27)
                           , QN => n136);
   Q_reg_26_inst : DFFR_X1 port map( D => n105, CK => CK, RN => n99, Q => Q(26)
                           , QN => n137);
   Q_reg_25_inst : DFFR_X1 port map( D => n106, CK => CK, RN => n99, Q => Q(25)
                           , QN => n138);
   Q_reg_24_inst : DFFR_X1 port map( D => n107, CK => CK, RN => n99, Q => Q(24)
                           , QN => n139);
   Q_reg_23_inst : DFFR_X1 port map( D => n108, CK => CK, RN => n98, Q => Q(23)
                           , QN => n140);
   Q_reg_22_inst : DFFR_X1 port map( D => n109, CK => CK, RN => n98, Q => Q(22)
                           , QN => n141);
   Q_reg_21_inst : DFFR_X1 port map( D => n110, CK => CK, RN => n98, Q => Q(21)
                           , QN => n142);
   Q_reg_20_inst : DFFR_X1 port map( D => n111, CK => CK, RN => n98, Q => Q(20)
                           , QN => n143);
   Q_reg_19_inst : DFFR_X1 port map( D => n112, CK => CK, RN => n98, Q => Q(19)
                           , QN => n144);
   Q_reg_18_inst : DFFR_X1 port map( D => n113, CK => CK, RN => n98, Q => Q(18)
                           , QN => n145);
   Q_reg_17_inst : DFFR_X1 port map( D => n114, CK => CK, RN => n98, Q => Q(17)
                           , QN => n146);
   Q_reg_16_inst : DFFR_X1 port map( D => n115, CK => CK, RN => n98, Q => Q(16)
                           , QN => n147);
   Q_reg_15_inst : DFFR_X1 port map( D => n116, CK => CK, RN => n98, Q => Q(15)
                           , QN => n148);
   Q_reg_14_inst : DFFR_X1 port map( D => n117, CK => CK, RN => n98, Q => Q(14)
                           , QN => n149);
   Q_reg_13_inst : DFFR_X1 port map( D => n118, CK => CK, RN => n98, Q => Q(13)
                           , QN => n150);
   Q_reg_12_inst : DFFR_X1 port map( D => n119, CK => CK, RN => n98, Q => Q(12)
                           , QN => n151);
   Q_reg_11_inst : DFFR_X1 port map( D => n120, CK => CK, RN => n97, Q => Q(11)
                           , QN => n152);
   Q_reg_10_inst : DFFR_X1 port map( D => n121, CK => CK, RN => n97, Q => Q(10)
                           , QN => n153);
   Q_reg_9_inst : DFFR_X1 port map( D => n122, CK => CK, RN => n97, Q => Q(9), 
                           QN => n154);
   Q_reg_8_inst : DFFR_X1 port map( D => n123, CK => CK, RN => n97, Q => Q(8), 
                           QN => n155);
   Q_reg_7_inst : DFFR_X1 port map( D => n124, CK => CK, RN => n97, Q => Q(7), 
                           QN => n156);
   Q_reg_6_inst : DFFR_X1 port map( D => n125, CK => CK, RN => n97, Q => Q(6), 
                           QN => n157);
   Q_reg_5_inst : DFFR_X1 port map( D => n126, CK => CK, RN => n97, Q => Q(5), 
                           QN => n158);
   Q_reg_4_inst : DFFR_X1 port map( D => n127, CK => CK, RN => n97, Q => Q(4), 
                           QN => n159);
   Q_reg_3_inst : DFFR_X1 port map( D => n128, CK => CK, RN => n97, Q => Q(3), 
                           QN => n160);
   Q_reg_2_inst : DFFR_X1 port map( D => n129, CK => CK, RN => n97, Q => Q(2), 
                           QN => n161);
   Q_reg_1_inst : DFFR_X1 port map( D => n130, CK => CK, RN => n97, Q => Q(1), 
                           QN => n162);
   Q_reg_0_inst : DFFR_X1 port map( D => n131, CK => CK, RN => n97, Q => Q(0), 
                           QN => n163);
   U2 : BUF_X1 port map( A => RESET, Z => n97);
   U3 : BUF_X1 port map( A => RESET, Z => n98);
   U4 : BUF_X1 port map( A => RESET, Z => n99);
   U5 : OAI21_X1 port map( B1 => n163, B2 => ENABLE, A => n195, ZN => n131);
   U6 : NAND2_X1 port map( A1 => ENABLE, A2 => D(0), ZN => n195);
   U7 : OAI21_X1 port map( B1 => n162, B2 => ENABLE, A => n194, ZN => n130);
   U8 : NAND2_X1 port map( A1 => D(1), A2 => ENABLE, ZN => n194);
   U9 : OAI21_X1 port map( B1 => n161, B2 => ENABLE, A => n193, ZN => n129);
   U10 : NAND2_X1 port map( A1 => D(2), A2 => ENABLE, ZN => n193);
   U11 : OAI21_X1 port map( B1 => n160, B2 => ENABLE, A => n192, ZN => n128);
   U12 : NAND2_X1 port map( A1 => D(3), A2 => ENABLE, ZN => n192);
   U13 : OAI21_X1 port map( B1 => n159, B2 => ENABLE, A => n191, ZN => n127);
   U14 : NAND2_X1 port map( A1 => D(4), A2 => ENABLE, ZN => n191);
   U15 : OAI21_X1 port map( B1 => n158, B2 => ENABLE, A => n190, ZN => n126);
   U16 : NAND2_X1 port map( A1 => D(5), A2 => ENABLE, ZN => n190);
   U17 : OAI21_X1 port map( B1 => n157, B2 => ENABLE, A => n189, ZN => n125);
   U18 : NAND2_X1 port map( A1 => D(6), A2 => ENABLE, ZN => n189);
   U19 : OAI21_X1 port map( B1 => n156, B2 => ENABLE, A => n188, ZN => n124);
   U20 : NAND2_X1 port map( A1 => D(7), A2 => ENABLE, ZN => n188);
   U21 : OAI21_X1 port map( B1 => n155, B2 => ENABLE, A => n187, ZN => n123);
   U22 : NAND2_X1 port map( A1 => D(8), A2 => ENABLE, ZN => n187);
   U23 : OAI21_X1 port map( B1 => n154, B2 => ENABLE, A => n186, ZN => n122);
   U24 : NAND2_X1 port map( A1 => D(9), A2 => ENABLE, ZN => n186);
   U25 : OAI21_X1 port map( B1 => n153, B2 => ENABLE, A => n185, ZN => n121);
   U26 : NAND2_X1 port map( A1 => D(10), A2 => ENABLE, ZN => n185);
   U27 : OAI21_X1 port map( B1 => n152, B2 => ENABLE, A => n184, ZN => n120);
   U28 : NAND2_X1 port map( A1 => D(11), A2 => ENABLE, ZN => n184);
   U29 : OAI21_X1 port map( B1 => n151, B2 => ENABLE, A => n183, ZN => n119);
   U30 : NAND2_X1 port map( A1 => D(12), A2 => ENABLE, ZN => n183);
   U31 : OAI21_X1 port map( B1 => n150, B2 => ENABLE, A => n182, ZN => n118);
   U32 : NAND2_X1 port map( A1 => D(13), A2 => ENABLE, ZN => n182);
   U33 : OAI21_X1 port map( B1 => n149, B2 => ENABLE, A => n181, ZN => n117);
   U34 : NAND2_X1 port map( A1 => D(14), A2 => ENABLE, ZN => n181);
   U35 : OAI21_X1 port map( B1 => n148, B2 => ENABLE, A => n180, ZN => n116);
   U36 : NAND2_X1 port map( A1 => D(15), A2 => ENABLE, ZN => n180);
   U37 : OAI21_X1 port map( B1 => n147, B2 => ENABLE, A => n179, ZN => n115);
   U38 : NAND2_X1 port map( A1 => D(16), A2 => ENABLE, ZN => n179);
   U39 : OAI21_X1 port map( B1 => n146, B2 => ENABLE, A => n178, ZN => n114);
   U40 : NAND2_X1 port map( A1 => D(17), A2 => ENABLE, ZN => n178);
   U41 : OAI21_X1 port map( B1 => n145, B2 => ENABLE, A => n177, ZN => n113);
   U42 : NAND2_X1 port map( A1 => D(18), A2 => ENABLE, ZN => n177);
   U43 : OAI21_X1 port map( B1 => n144, B2 => ENABLE, A => n176, ZN => n112);
   U44 : NAND2_X1 port map( A1 => D(19), A2 => ENABLE, ZN => n176);
   U45 : OAI21_X1 port map( B1 => n143, B2 => ENABLE, A => n175, ZN => n111);
   U46 : NAND2_X1 port map( A1 => D(20), A2 => ENABLE, ZN => n175);
   U47 : OAI21_X1 port map( B1 => n142, B2 => ENABLE, A => n174, ZN => n110);
   U48 : NAND2_X1 port map( A1 => D(21), A2 => ENABLE, ZN => n174);
   U49 : OAI21_X1 port map( B1 => n141, B2 => ENABLE, A => n173, ZN => n109);
   U50 : NAND2_X1 port map( A1 => D(22), A2 => ENABLE, ZN => n173);
   U51 : OAI21_X1 port map( B1 => n140, B2 => ENABLE, A => n172, ZN => n108);
   U52 : NAND2_X1 port map( A1 => D(23), A2 => ENABLE, ZN => n172);
   U53 : OAI21_X1 port map( B1 => n139, B2 => ENABLE, A => n171, ZN => n107);
   U54 : NAND2_X1 port map( A1 => D(24), A2 => ENABLE, ZN => n171);
   U55 : OAI21_X1 port map( B1 => n138, B2 => ENABLE, A => n170, ZN => n106);
   U56 : NAND2_X1 port map( A1 => D(25), A2 => ENABLE, ZN => n170);
   U57 : OAI21_X1 port map( B1 => n137, B2 => ENABLE, A => n169, ZN => n105);
   U58 : NAND2_X1 port map( A1 => D(26), A2 => ENABLE, ZN => n169);
   U59 : OAI21_X1 port map( B1 => n136, B2 => ENABLE, A => n168, ZN => n104);
   U60 : NAND2_X1 port map( A1 => D(27), A2 => ENABLE, ZN => n168);
   U61 : OAI21_X1 port map( B1 => n135, B2 => ENABLE, A => n167, ZN => n103);
   U62 : NAND2_X1 port map( A1 => D(28), A2 => ENABLE, ZN => n167);
   U63 : OAI21_X1 port map( B1 => n134, B2 => ENABLE, A => n166, ZN => n102);
   U64 : NAND2_X1 port map( A1 => D(29), A2 => ENABLE, ZN => n166);
   U65 : OAI21_X1 port map( B1 => n133, B2 => ENABLE, A => n165, ZN => n101);
   U66 : NAND2_X1 port map( A1 => D(30), A2 => ENABLE, ZN => n165);
   U67 : OAI21_X1 port map( B1 => n132, B2 => ENABLE, A => n164, ZN => n100);
   U68 : NAND2_X1 port map( A1 => D(31), A2 => ENABLE, ZN => n164);

end SYN_ASYNCHBEHAV;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity regFFD_NBIT32_1 is

   port( CK, RESET, ENABLE : in std_logic;  D : in std_logic_vector (31 downto 
         0);  Q : out std_logic_vector (31 downto 0));

end regFFD_NBIT32_1;

architecture SYN_ASYNCHBEHAV of regFFD_NBIT32_1 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, 
      n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, 
      n121, n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, 
      n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, 
      n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, 
      n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, 
      n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, 
      n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, 
      n193, n194, n195 : std_logic;

begin
   
   Q_reg_31_inst : DFFR_X1 port map( D => n100, CK => CK, RN => n99, Q => Q(31)
                           , QN => n132);
   Q_reg_30_inst : DFFR_X1 port map( D => n101, CK => CK, RN => n99, Q => Q(30)
                           , QN => n133);
   Q_reg_29_inst : DFFR_X1 port map( D => n102, CK => CK, RN => n99, Q => Q(29)
                           , QN => n134);
   Q_reg_28_inst : DFFR_X1 port map( D => n103, CK => CK, RN => n99, Q => Q(28)
                           , QN => n135);
   Q_reg_27_inst : DFFR_X1 port map( D => n104, CK => CK, RN => n99, Q => Q(27)
                           , QN => n136);
   Q_reg_26_inst : DFFR_X1 port map( D => n105, CK => CK, RN => n99, Q => Q(26)
                           , QN => n137);
   Q_reg_25_inst : DFFR_X1 port map( D => n106, CK => CK, RN => n99, Q => Q(25)
                           , QN => n138);
   Q_reg_24_inst : DFFR_X1 port map( D => n107, CK => CK, RN => n99, Q => Q(24)
                           , QN => n139);
   Q_reg_23_inst : DFFR_X1 port map( D => n108, CK => CK, RN => n98, Q => Q(23)
                           , QN => n140);
   Q_reg_22_inst : DFFR_X1 port map( D => n109, CK => CK, RN => n98, Q => Q(22)
                           , QN => n141);
   Q_reg_21_inst : DFFR_X1 port map( D => n110, CK => CK, RN => n98, Q => Q(21)
                           , QN => n142);
   Q_reg_20_inst : DFFR_X1 port map( D => n111, CK => CK, RN => n98, Q => Q(20)
                           , QN => n143);
   Q_reg_19_inst : DFFR_X1 port map( D => n112, CK => CK, RN => n98, Q => Q(19)
                           , QN => n144);
   Q_reg_18_inst : DFFR_X1 port map( D => n113, CK => CK, RN => n98, Q => Q(18)
                           , QN => n145);
   Q_reg_17_inst : DFFR_X1 port map( D => n114, CK => CK, RN => n98, Q => Q(17)
                           , QN => n146);
   Q_reg_16_inst : DFFR_X1 port map( D => n115, CK => CK, RN => n98, Q => Q(16)
                           , QN => n147);
   Q_reg_15_inst : DFFR_X1 port map( D => n116, CK => CK, RN => n98, Q => Q(15)
                           , QN => n148);
   Q_reg_14_inst : DFFR_X1 port map( D => n117, CK => CK, RN => n98, Q => Q(14)
                           , QN => n149);
   Q_reg_13_inst : DFFR_X1 port map( D => n118, CK => CK, RN => n98, Q => Q(13)
                           , QN => n150);
   Q_reg_12_inst : DFFR_X1 port map( D => n119, CK => CK, RN => n98, Q => Q(12)
                           , QN => n151);
   Q_reg_11_inst : DFFR_X1 port map( D => n120, CK => CK, RN => n97, Q => Q(11)
                           , QN => n152);
   Q_reg_10_inst : DFFR_X1 port map( D => n121, CK => CK, RN => n97, Q => Q(10)
                           , QN => n153);
   Q_reg_9_inst : DFFR_X1 port map( D => n122, CK => CK, RN => n97, Q => Q(9), 
                           QN => n154);
   Q_reg_8_inst : DFFR_X1 port map( D => n123, CK => CK, RN => n97, Q => Q(8), 
                           QN => n155);
   Q_reg_7_inst : DFFR_X1 port map( D => n124, CK => CK, RN => n97, Q => Q(7), 
                           QN => n156);
   Q_reg_6_inst : DFFR_X1 port map( D => n125, CK => CK, RN => n97, Q => Q(6), 
                           QN => n157);
   Q_reg_5_inst : DFFR_X1 port map( D => n126, CK => CK, RN => n97, Q => Q(5), 
                           QN => n158);
   Q_reg_4_inst : DFFR_X1 port map( D => n127, CK => CK, RN => n97, Q => Q(4), 
                           QN => n159);
   Q_reg_3_inst : DFFR_X1 port map( D => n128, CK => CK, RN => n97, Q => Q(3), 
                           QN => n160);
   Q_reg_2_inst : DFFR_X1 port map( D => n129, CK => CK, RN => n97, Q => Q(2), 
                           QN => n161);
   Q_reg_1_inst : DFFR_X1 port map( D => n130, CK => CK, RN => n97, Q => Q(1), 
                           QN => n162);
   Q_reg_0_inst : DFFR_X1 port map( D => n131, CK => CK, RN => n97, Q => Q(0), 
                           QN => n163);
   U2 : BUF_X1 port map( A => RESET, Z => n97);
   U3 : BUF_X1 port map( A => RESET, Z => n98);
   U4 : BUF_X1 port map( A => RESET, Z => n99);
   U5 : OAI21_X1 port map( B1 => n163, B2 => ENABLE, A => n195, ZN => n131);
   U6 : NAND2_X1 port map( A1 => ENABLE, A2 => D(0), ZN => n195);
   U7 : OAI21_X1 port map( B1 => n162, B2 => ENABLE, A => n194, ZN => n130);
   U8 : NAND2_X1 port map( A1 => D(1), A2 => ENABLE, ZN => n194);
   U9 : OAI21_X1 port map( B1 => n161, B2 => ENABLE, A => n193, ZN => n129);
   U10 : NAND2_X1 port map( A1 => D(2), A2 => ENABLE, ZN => n193);
   U11 : OAI21_X1 port map( B1 => n160, B2 => ENABLE, A => n192, ZN => n128);
   U12 : NAND2_X1 port map( A1 => D(3), A2 => ENABLE, ZN => n192);
   U13 : OAI21_X1 port map( B1 => n159, B2 => ENABLE, A => n191, ZN => n127);
   U14 : NAND2_X1 port map( A1 => D(4), A2 => ENABLE, ZN => n191);
   U15 : OAI21_X1 port map( B1 => n158, B2 => ENABLE, A => n190, ZN => n126);
   U16 : NAND2_X1 port map( A1 => D(5), A2 => ENABLE, ZN => n190);
   U17 : OAI21_X1 port map( B1 => n157, B2 => ENABLE, A => n189, ZN => n125);
   U18 : NAND2_X1 port map( A1 => D(6), A2 => ENABLE, ZN => n189);
   U19 : OAI21_X1 port map( B1 => n156, B2 => ENABLE, A => n188, ZN => n124);
   U20 : NAND2_X1 port map( A1 => D(7), A2 => ENABLE, ZN => n188);
   U21 : OAI21_X1 port map( B1 => n155, B2 => ENABLE, A => n187, ZN => n123);
   U22 : NAND2_X1 port map( A1 => D(8), A2 => ENABLE, ZN => n187);
   U23 : OAI21_X1 port map( B1 => n154, B2 => ENABLE, A => n186, ZN => n122);
   U24 : NAND2_X1 port map( A1 => D(9), A2 => ENABLE, ZN => n186);
   U25 : OAI21_X1 port map( B1 => n153, B2 => ENABLE, A => n185, ZN => n121);
   U26 : NAND2_X1 port map( A1 => D(10), A2 => ENABLE, ZN => n185);
   U27 : OAI21_X1 port map( B1 => n152, B2 => ENABLE, A => n184, ZN => n120);
   U28 : NAND2_X1 port map( A1 => D(11), A2 => ENABLE, ZN => n184);
   U29 : OAI21_X1 port map( B1 => n151, B2 => ENABLE, A => n183, ZN => n119);
   U30 : NAND2_X1 port map( A1 => D(12), A2 => ENABLE, ZN => n183);
   U31 : OAI21_X1 port map( B1 => n150, B2 => ENABLE, A => n182, ZN => n118);
   U32 : NAND2_X1 port map( A1 => D(13), A2 => ENABLE, ZN => n182);
   U33 : OAI21_X1 port map( B1 => n149, B2 => ENABLE, A => n181, ZN => n117);
   U34 : NAND2_X1 port map( A1 => D(14), A2 => ENABLE, ZN => n181);
   U35 : OAI21_X1 port map( B1 => n148, B2 => ENABLE, A => n180, ZN => n116);
   U36 : NAND2_X1 port map( A1 => D(15), A2 => ENABLE, ZN => n180);
   U37 : OAI21_X1 port map( B1 => n147, B2 => ENABLE, A => n179, ZN => n115);
   U38 : NAND2_X1 port map( A1 => D(16), A2 => ENABLE, ZN => n179);
   U39 : OAI21_X1 port map( B1 => n146, B2 => ENABLE, A => n178, ZN => n114);
   U40 : NAND2_X1 port map( A1 => D(17), A2 => ENABLE, ZN => n178);
   U41 : OAI21_X1 port map( B1 => n145, B2 => ENABLE, A => n177, ZN => n113);
   U42 : NAND2_X1 port map( A1 => D(18), A2 => ENABLE, ZN => n177);
   U43 : OAI21_X1 port map( B1 => n144, B2 => ENABLE, A => n176, ZN => n112);
   U44 : NAND2_X1 port map( A1 => D(19), A2 => ENABLE, ZN => n176);
   U45 : OAI21_X1 port map( B1 => n143, B2 => ENABLE, A => n175, ZN => n111);
   U46 : NAND2_X1 port map( A1 => D(20), A2 => ENABLE, ZN => n175);
   U47 : OAI21_X1 port map( B1 => n142, B2 => ENABLE, A => n174, ZN => n110);
   U48 : NAND2_X1 port map( A1 => D(21), A2 => ENABLE, ZN => n174);
   U49 : OAI21_X1 port map( B1 => n141, B2 => ENABLE, A => n173, ZN => n109);
   U50 : NAND2_X1 port map( A1 => D(22), A2 => ENABLE, ZN => n173);
   U51 : OAI21_X1 port map( B1 => n140, B2 => ENABLE, A => n172, ZN => n108);
   U52 : NAND2_X1 port map( A1 => D(23), A2 => ENABLE, ZN => n172);
   U53 : OAI21_X1 port map( B1 => n139, B2 => ENABLE, A => n171, ZN => n107);
   U54 : NAND2_X1 port map( A1 => D(24), A2 => ENABLE, ZN => n171);
   U55 : OAI21_X1 port map( B1 => n138, B2 => ENABLE, A => n170, ZN => n106);
   U56 : NAND2_X1 port map( A1 => D(25), A2 => ENABLE, ZN => n170);
   U57 : OAI21_X1 port map( B1 => n137, B2 => ENABLE, A => n169, ZN => n105);
   U58 : NAND2_X1 port map( A1 => D(26), A2 => ENABLE, ZN => n169);
   U59 : OAI21_X1 port map( B1 => n136, B2 => ENABLE, A => n168, ZN => n104);
   U60 : NAND2_X1 port map( A1 => D(27), A2 => ENABLE, ZN => n168);
   U61 : OAI21_X1 port map( B1 => n135, B2 => ENABLE, A => n167, ZN => n103);
   U62 : NAND2_X1 port map( A1 => D(28), A2 => ENABLE, ZN => n167);
   U63 : OAI21_X1 port map( B1 => n134, B2 => ENABLE, A => n166, ZN => n102);
   U64 : NAND2_X1 port map( A1 => D(29), A2 => ENABLE, ZN => n166);
   U65 : OAI21_X1 port map( B1 => n133, B2 => ENABLE, A => n165, ZN => n101);
   U66 : NAND2_X1 port map( A1 => D(30), A2 => ENABLE, ZN => n165);
   U67 : OAI21_X1 port map( B1 => n132, B2 => ENABLE, A => n164, ZN => n100);
   U68 : NAND2_X1 port map( A1 => D(31), A2 => ENABLE, ZN => n164);

end SYN_ASYNCHBEHAV;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_GENERIC_NBIT4_0 is

   port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (3 downto 0));

end MUX21_GENERIC_NBIT4_0;

architecture SYN_struct of MUX21_GENERIC_NBIT4_0 is

   component MUX21_29
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_30
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_31
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_32
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;

begin
   
   gen1_0 : MUX21_32 port map( A => A(0), B => B(0), S => SEL, Y => Y(0));
   gen1_1 : MUX21_31 port map( A => A(1), B => B(1), S => SEL, Y => Y(1));
   gen1_2 : MUX21_30 port map( A => A(2), B => B(2), S => SEL, Y => Y(2));
   gen1_3 : MUX21_29 port map( A => A(3), B => B(3), S => SEL, Y => Y(3));

end SYN_struct;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity RCA_NBIT4_0 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_NBIT4_0;

architecture SYN_BEHAVIORAL of RCA_NBIT4_0 is

   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal add_1_root_add_52_2_carry_1_port, add_1_root_add_52_2_carry_2_port, 
      add_1_root_add_52_2_carry_3_port : std_logic;

begin
   
   add_1_root_add_52_2_U1_0 : FA_X1 port map( A => A(0), B => B(0), CI => Ci, 
                           CO => add_1_root_add_52_2_carry_1_port, S => S(0));
   add_1_root_add_52_2_U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => 
                           add_1_root_add_52_2_carry_1_port, CO => 
                           add_1_root_add_52_2_carry_2_port, S => S(1));
   add_1_root_add_52_2_U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => 
                           add_1_root_add_52_2_carry_2_port, CO => 
                           add_1_root_add_52_2_carry_3_port, S => S(2));
   add_1_root_add_52_2_U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => 
                           add_1_root_add_52_2_carry_3_port, CO => Co, S => 
                           S(3));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity P_0 is

   port( p1, P2 : in std_logic;  Co : out std_logic);

end P_0;

architecture SYN_behave of P_0 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => p1, A2 => P2, ZN => Co);

end SYN_behave;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity CSB_NBIT4_0 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0));

end CSB_NBIT4_0;

architecture SYN_STRUCTURAL of CSB_NBIT4_0 is

   component MUX21_GENERIC_NBIT4_0
      port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component RCA_NBIT4_15
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCA_NBIT4_0
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, out_rca0_3_port, out_rca0_2_port, 
      out_rca0_1_port, out_rca0_0_port, out_rca1_3_port, out_rca1_2_port, 
      out_rca1_1_port, out_rca1_0_port, n_1041, n_1042 : std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA0 : RCA_NBIT4_0 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), A(0) 
                           => A(0), B(3) => B(3), B(2) => B(2), B(1) => B(1), 
                           B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           out_rca0_3_port, S(2) => out_rca0_2_port, S(1) => 
                           out_rca0_1_port, S(0) => out_rca0_0_port, Co => 
                           n_1041);
   RCA1 : RCA_NBIT4_15 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), A(0)
                           => A(0), B(3) => B(3), B(2) => B(2), B(1) => B(1), 
                           B(0) => B(0), Ci => X_Logic1_port, S(3) => 
                           out_rca1_3_port, S(2) => out_rca1_2_port, S(1) => 
                           out_rca1_1_port, S(0) => out_rca1_0_port, Co => 
                           n_1042);
   MUXCin : MUX21_GENERIC_NBIT4_0 port map( A(3) => out_rca1_3_port, A(2) => 
                           out_rca1_2_port, A(1) => out_rca1_1_port, A(0) => 
                           out_rca1_0_port, B(3) => out_rca0_3_port, B(2) => 
                           out_rca0_2_port, B(1) => out_rca0_1_port, B(0) => 
                           out_rca0_0_port, SEL => Ci, Y(3) => S(3), Y(2) => 
                           S(2), Y(1) => S(1), Y(0) => S(0));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity PG_0 is

   port( G1, P1, G2, P2 : in std_logic;  gout, pout : out std_logic);

end PG_0;

architecture SYN_arch of PG_0 is

   component P_0
      port( p1, P2 : in std_logic;  Co : out std_logic);
   end component;
   
   component G_43
      port( G1, P, G2 : in std_logic;  Co : out std_logic);
   end component;

begin
   
   g_comp : G_43 port map( G1 => G1, P => P1, G2 => G2, Co => gout);
   p_comp : P_0 port map( p1 => P1, P2 => P2, Co => pout);

end SYN_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity G_0 is

   port( G1, P, G2 : in std_logic;  Co : out std_logic);

end G_0;

architecture SYN_behave of G_0 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n2, ZN => Co);
   U2 : AOI21_X1 port map( B1 => P, B2 => G2, A => G1, ZN => n2);

end SYN_behave;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity SUM_GENERATOR_NBIT_PER_BLOCK4_NBLOCKS8 is

   port( A, B : in std_logic_vector (31 downto 0);  Ci : in std_logic_vector (7
         downto 0);  S : out std_logic_vector (31 downto 0));

end SUM_GENERATOR_NBIT_PER_BLOCK4_NBLOCKS8;

architecture SYN_STRUCTURAL of SUM_GENERATOR_NBIT_PER_BLOCK4_NBLOCKS8 is

   component CSB_NBIT4_1
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component CSB_NBIT4_2
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component CSB_NBIT4_3
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component CSB_NBIT4_4
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component CSB_NBIT4_5
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component CSB_NBIT4_6
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component CSB_NBIT4_7
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component CSB_NBIT4_0
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0));
   end component;

begin
   
   CSBI_0 : CSB_NBIT4_0 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => Ci(0), S(3) => S(3), S(2) 
                           => S(2), S(1) => S(1), S(0) => S(0));
   CSBI_1 : CSB_NBIT4_7 port map( A(3) => A(7), A(2) => A(6), A(1) => A(5), 
                           A(0) => A(4), B(3) => B(7), B(2) => B(6), B(1) => 
                           B(5), B(0) => B(4), Ci => Ci(1), S(3) => S(7), S(2) 
                           => S(6), S(1) => S(5), S(0) => S(4));
   CSBI_2 : CSB_NBIT4_6 port map( A(3) => A(11), A(2) => A(10), A(1) => A(9), 
                           A(0) => A(8), B(3) => B(11), B(2) => B(10), B(1) => 
                           B(9), B(0) => B(8), Ci => Ci(2), S(3) => S(11), S(2)
                           => S(10), S(1) => S(9), S(0) => S(8));
   CSBI_3 : CSB_NBIT4_5 port map( A(3) => A(15), A(2) => A(14), A(1) => A(13), 
                           A(0) => A(12), B(3) => B(15), B(2) => B(14), B(1) =>
                           B(13), B(0) => B(12), Ci => Ci(3), S(3) => S(15), 
                           S(2) => S(14), S(1) => S(13), S(0) => S(12));
   CSBI_4 : CSB_NBIT4_4 port map( A(3) => A(19), A(2) => A(18), A(1) => A(17), 
                           A(0) => A(16), B(3) => B(19), B(2) => B(18), B(1) =>
                           B(17), B(0) => B(16), Ci => Ci(4), S(3) => S(19), 
                           S(2) => S(18), S(1) => S(17), S(0) => S(16));
   CSBI_5 : CSB_NBIT4_3 port map( A(3) => A(23), A(2) => A(22), A(1) => A(21), 
                           A(0) => A(20), B(3) => B(23), B(2) => B(22), B(1) =>
                           B(21), B(0) => B(20), Ci => Ci(5), S(3) => S(23), 
                           S(2) => S(22), S(1) => S(21), S(0) => S(20));
   CSBI_6 : CSB_NBIT4_2 port map( A(3) => A(27), A(2) => A(26), A(1) => A(25), 
                           A(0) => A(24), B(3) => B(27), B(2) => B(26), B(1) =>
                           B(25), B(0) => B(24), Ci => Ci(6), S(3) => S(27), 
                           S(2) => S(26), S(1) => S(25), S(0) => S(24));
   CSBI_7 : CSB_NBIT4_1 port map( A(3) => A(31), A(2) => A(30), A(1) => A(29), 
                           A(0) => A(28), B(3) => B(31), B(2) => B(30), B(1) =>
                           B(29), B(0) => B(28), Ci => Ci(7), S(3) => S(31), 
                           S(2) => S(30), S(1) => S(29), S(0) => S(28));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity CARRY_GENERATOR_NBIT32_NBIT_PER_BLOCK4 is

   port( A, B : in std_logic_vector (31 downto 0);  Cin : in std_logic;  Co : 
         out std_logic_vector (7 downto 0));

end CARRY_GENERATOR_NBIT32_NBIT_PER_BLOCK4;

architecture SYN_arch of CARRY_GENERATOR_NBIT32_NBIT_PER_BLOCK4 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component G_44
      port( G1, P, G2 : in std_logic;  Co : out std_logic);
   end component;
   
   component G_45
      port( G1, P, G2 : in std_logic;  Co : out std_logic);
   end component;
   
   component G_46
      port( G1, P, G2 : in std_logic;  Co : out std_logic);
   end component;
   
   component G_47
      port( G1, P, G2 : in std_logic;  Co : out std_logic);
   end component;
   
   component PG_1
      port( G1, P1, G2, P2 : in std_logic;  gout, pout : out std_logic);
   end component;
   
   component PG_2
      port( G1, P1, G2, P2 : in std_logic;  gout, pout : out std_logic);
   end component;
   
   component G_48
      port( G1, P, G2 : in std_logic;  Co : out std_logic);
   end component;
   
   component G_49
      port( G1, P, G2 : in std_logic;  Co : out std_logic);
   end component;
   
   component PG_3
      port( G1, P1, G2, P2 : in std_logic;  gout, pout : out std_logic);
   end component;
   
   component PG_4
      port( G1, P1, G2, P2 : in std_logic;  gout, pout : out std_logic);
   end component;
   
   component PG_5
      port( G1, P1, G2, P2 : in std_logic;  gout, pout : out std_logic);
   end component;
   
   component G_50
      port( G1, P, G2 : in std_logic;  Co : out std_logic);
   end component;
   
   component PG_6
      port( G1, P1, G2, P2 : in std_logic;  gout, pout : out std_logic);
   end component;
   
   component PG_7
      port( G1, P1, G2, P2 : in std_logic;  gout, pout : out std_logic);
   end component;
   
   component PG_8
      port( G1, P1, G2, P2 : in std_logic;  gout, pout : out std_logic);
   end component;
   
   component PG_9
      port( G1, P1, G2, P2 : in std_logic;  gout, pout : out std_logic);
   end component;
   
   component PG_10
      port( G1, P1, G2, P2 : in std_logic;  gout, pout : out std_logic);
   end component;
   
   component PG_11
      port( G1, P1, G2, P2 : in std_logic;  gout, pout : out std_logic);
   end component;
   
   component PG_12
      port( G1, P1, G2, P2 : in std_logic;  gout, pout : out std_logic);
   end component;
   
   component G_51
      port( G1, P, G2 : in std_logic;  Co : out std_logic);
   end component;
   
   component PG_13
      port( G1, P1, G2, P2 : in std_logic;  gout, pout : out std_logic);
   end component;
   
   component PG_14
      port( G1, P1, G2, P2 : in std_logic;  gout, pout : out std_logic);
   end component;
   
   component PG_15
      port( G1, P1, G2, P2 : in std_logic;  gout, pout : out std_logic);
   end component;
   
   component PG_16
      port( G1, P1, G2, P2 : in std_logic;  gout, pout : out std_logic);
   end component;
   
   component PG_17
      port( G1, P1, G2, P2 : in std_logic;  gout, pout : out std_logic);
   end component;
   
   component PG_18
      port( G1, P1, G2, P2 : in std_logic;  gout, pout : out std_logic);
   end component;
   
   component PG_19
      port( G1, P1, G2, P2 : in std_logic;  gout, pout : out std_logic);
   end component;
   
   component PG_20
      port( G1, P1, G2, P2 : in std_logic;  gout, pout : out std_logic);
   end component;
   
   component PG_21
      port( G1, P1, G2, P2 : in std_logic;  gout, pout : out std_logic);
   end component;
   
   component PG_22
      port( G1, P1, G2, P2 : in std_logic;  gout, pout : out std_logic);
   end component;
   
   component PG_23
      port( G1, P1, G2, P2 : in std_logic;  gout, pout : out std_logic);
   end component;
   
   component PG_24
      port( G1, P1, G2, P2 : in std_logic;  gout, pout : out std_logic);
   end component;
   
   component PG_25
      port( G1, P1, G2, P2 : in std_logic;  gout, pout : out std_logic);
   end component;
   
   component PG_26
      port( G1, P1, G2, P2 : in std_logic;  gout, pout : out std_logic);
   end component;
   
   component PG_27
      port( G1, P1, G2, P2 : in std_logic;  gout, pout : out std_logic);
   end component;
   
   component PG_28
      port( G1, P1, G2, P2 : in std_logic;  gout, pout : out std_logic);
   end component;
   
   component PG_29
      port( G1, P1, G2, P2 : in std_logic;  gout, pout : out std_logic);
   end component;
   
   component PG_30
      port( G1, P1, G2, P2 : in std_logic;  gout, pout : out std_logic);
   end component;
   
   component PG_31
      port( G1, P1, G2, P2 : in std_logic;  gout, pout : out std_logic);
   end component;
   
   component PG_32
      port( G1, P1, G2, P2 : in std_logic;  gout, pout : out std_logic);
   end component;
   
   component PG_33
      port( G1, P1, G2, P2 : in std_logic;  gout, pout : out std_logic);
   end component;
   
   component PG_34
      port( G1, P1, G2, P2 : in std_logic;  gout, pout : out std_logic);
   end component;
   
   component PG_35
      port( G1, P1, G2, P2 : in std_logic;  gout, pout : out std_logic);
   end component;
   
   component PG_36
      port( G1, P1, G2, P2 : in std_logic;  gout, pout : out std_logic);
   end component;
   
   component PG_37
      port( G1, P1, G2, P2 : in std_logic;  gout, pout : out std_logic);
   end component;
   
   component PG_38
      port( G1, P1, G2, P2 : in std_logic;  gout, pout : out std_logic);
   end component;
   
   component PG_39
      port( G1, P1, G2, P2 : in std_logic;  gout, pout : out std_logic);
   end component;
   
   component PG_40
      port( G1, P1, G2, P2 : in std_logic;  gout, pout : out std_logic);
   end component;
   
   component PG_41
      port( G1, P1, G2, P2 : in std_logic;  gout, pout : out std_logic);
   end component;
   
   component PG_42
      port( G1, P1, G2, P2 : in std_logic;  gout, pout : out std_logic);
   end component;
   
   component G_52
      port( G1, P, G2 : in std_logic;  Co : out std_logic);
   end component;
   
   component PG_0
      port( G1, P1, G2, P2 : in std_logic;  gout, pout : out std_logic);
   end component;
   
   component G_0
      port( G1, P, G2 : in std_logic;  Co : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal X_Logic0_port, Co_7_port, Co_6_port, Co_5_port, Co_4_port, Co_3_port,
      Co_2_port, Co_1_port, Co_0_port, gi_32_4_port, gi_32_3_port, gi_32_2_port
      , gi_32_1_port, gi_32_0_port, gi_31_0_port, gi_30_0_port, gi_29_0_port, 
      gi_28_4_port, gi_28_2_port, gi_28_1_port, gi_28_0_port, gi_27_0_port, 
      gi_26_0_port, gi_25_0_port, gi_24_3_port, gi_24_2_port, gi_24_1_port, 
      gi_24_0_port, gi_23_0_port, gi_22_0_port, gi_21_0_port, gi_20_2_port, 
      gi_20_1_port, gi_20_0_port, gi_19_0_port, gi_18_0_port, gi_17_0_port, 
      gi_16_3_port, gi_16_2_port, gi_16_1_port, gi_16_0_port, gi_15_0_port, 
      gi_14_0_port, gi_13_0_port, gi_12_2_port, gi_12_1_port, gi_12_0_port, 
      gi_11_0_port, gi_10_0_port, gi_9_0_port, gi_8_2_port, gi_8_1_port, 
      gi_8_0_port, gi_7_0_port, gi_6_0_port, gi_5_0_port, gi_4_1_port, 
      gi_4_0_port, gi_3_0_port, gi_2_1_port, gi_2_0_port, gi_1_0_port, 
      gi_0_0_port, pi_32_4_port, pi_32_3_port, pi_32_2_port, pi_32_1_port, 
      pi_32_0_port, pi_31_0_port, pi_30_0_port, pi_29_0_port, pi_28_4_port, 
      pi_28_2_port, pi_28_1_port, pi_28_0_port, pi_27_0_port, pi_26_0_port, 
      pi_25_0_port, pi_24_3_port, pi_24_2_port, pi_24_1_port, pi_24_0_port, 
      pi_23_0_port, pi_22_0_port, pi_21_0_port, pi_20_2_port, pi_20_1_port, 
      pi_20_0_port, pi_19_0_port, pi_18_0_port, pi_17_0_port, pi_16_3_port, 
      pi_16_2_port, pi_16_1_port, pi_16_0_port, pi_15_0_port, pi_14_0_port, 
      pi_13_0_port, pi_12_2_port, pi_12_1_port, pi_12_0_port, pi_11_0_port, 
      pi_10_0_port, pi_9_0_port, pi_8_2_port, pi_8_1_port, pi_8_0_port, 
      pi_7_0_port, pi_6_0_port, pi_5_0_port, pi_4_1_port, pi_4_0_port, 
      pi_3_0_port, pi_2_0_port, pi_0_0_port, n_1043, n_1044, n_1045, n_1046, 
      n_1047, n_1048, n_1049, n_1050, n_1051, n_1052, n_1053, n_1054, n_1055, 
      n_1056, n_1057, n_1058, n_1059, n_1060, n_1061, n_1062, n_1063, n_1064, 
      n_1065, n_1066, n_1067, n_1068, n_1069, n_1070, n_1071, n_1072, n_1073, 
      n_1074, n_1075, n_1076, n_1077, n_1078, n_1079, n_1080, n_1081, n_1082, 
      n_1083, n_1084, n_1085, n_1086, n_1087, n_1088 : std_logic;

begin
   Co <= ( Co_7_port, Co_6_port, Co_5_port, Co_4_port, Co_3_port, Co_2_port, 
      Co_1_port, Co_0_port );
   
   X_Logic0_port <= '0';
   U34 : XOR2_X1 port map( A => B(8), B => A(8), Z => pi_9_0_port);
   U35 : XOR2_X1 port map( A => B(7), B => A(7), Z => pi_8_0_port);
   U36 : XOR2_X1 port map( A => B(6), B => A(6), Z => pi_7_0_port);
   U37 : XOR2_X1 port map( A => B(5), B => A(5), Z => pi_6_0_port);
   U38 : XOR2_X1 port map( A => B(4), B => A(4), Z => pi_5_0_port);
   U39 : XOR2_X1 port map( A => B(3), B => A(3), Z => pi_4_0_port);
   U40 : XOR2_X1 port map( A => B(2), B => A(2), Z => pi_3_0_port);
   U41 : XOR2_X1 port map( A => B(31), B => A(31), Z => pi_32_0_port);
   U42 : XOR2_X1 port map( A => B(30), B => A(30), Z => pi_31_0_port);
   U43 : XOR2_X1 port map( A => B(29), B => A(29), Z => pi_30_0_port);
   U44 : XOR2_X1 port map( A => B(1), B => A(1), Z => pi_2_0_port);
   U45 : XOR2_X1 port map( A => B(28), B => A(28), Z => pi_29_0_port);
   U46 : XOR2_X1 port map( A => B(27), B => A(27), Z => pi_28_0_port);
   U47 : XOR2_X1 port map( A => B(26), B => A(26), Z => pi_27_0_port);
   U48 : XOR2_X1 port map( A => B(25), B => A(25), Z => pi_26_0_port);
   U49 : XOR2_X1 port map( A => B(24), B => A(24), Z => pi_25_0_port);
   U50 : XOR2_X1 port map( A => B(23), B => A(23), Z => pi_24_0_port);
   U51 : XOR2_X1 port map( A => B(22), B => A(22), Z => pi_23_0_port);
   U52 : XOR2_X1 port map( A => B(21), B => A(21), Z => pi_22_0_port);
   U53 : XOR2_X1 port map( A => B(20), B => A(20), Z => pi_21_0_port);
   U54 : XOR2_X1 port map( A => B(19), B => A(19), Z => pi_20_0_port);
   U55 : XOR2_X1 port map( A => B(18), B => A(18), Z => pi_19_0_port);
   U56 : XOR2_X1 port map( A => B(17), B => A(17), Z => pi_18_0_port);
   U57 : XOR2_X1 port map( A => B(16), B => A(16), Z => pi_17_0_port);
   U58 : XOR2_X1 port map( A => B(15), B => A(15), Z => pi_16_0_port);
   U59 : XOR2_X1 port map( A => B(14), B => A(14), Z => pi_15_0_port);
   U60 : XOR2_X1 port map( A => B(13), B => A(13), Z => pi_14_0_port);
   U61 : XOR2_X1 port map( A => B(12), B => A(12), Z => pi_13_0_port);
   U62 : XOR2_X1 port map( A => B(11), B => A(11), Z => pi_12_0_port);
   U63 : XOR2_X1 port map( A => B(10), B => A(10), Z => pi_11_0_port);
   U64 : XOR2_X1 port map( A => B(9), B => A(9), Z => pi_10_0_port);
   U65 : XOR2_X1 port map( A => B(0), B => A(0), Z => pi_0_0_port);
   g_port0_0_1 : G_0 port map( G1 => gi_0_0_port, P => pi_0_0_port, G2 => Cin, 
                           Co => gi_1_0_port);
   pg_port2_1_1 : PG_0 port map( G1 => gi_1_0_port, P1 => X_Logic0_port, G2 => 
                           gi_0_0_port, P2 => pi_0_0_port, gout => n_1043, pout
                           => n_1044);
   g_port1_1_2 : G_52 port map( G1 => gi_2_0_port, P => pi_2_0_port, G2 => 
                           gi_1_0_port, Co => gi_2_1_port);
   pg_port2_1_3 : PG_42 port map( G1 => gi_3_0_port, P1 => pi_3_0_port, G2 => 
                           gi_2_0_port, P2 => pi_2_0_port, gout => n_1045, pout
                           => n_1046);
   pg_port2_1_4 : PG_41 port map( G1 => gi_4_0_port, P1 => pi_4_0_port, G2 => 
                           gi_3_0_port, P2 => pi_3_0_port, gout => gi_4_1_port,
                           pout => pi_4_1_port);
   pg_port2_1_5 : PG_40 port map( G1 => gi_5_0_port, P1 => pi_5_0_port, G2 => 
                           gi_4_0_port, P2 => pi_4_0_port, gout => n_1047, pout
                           => n_1048);
   pg_port2_1_6 : PG_39 port map( G1 => gi_6_0_port, P1 => pi_6_0_port, G2 => 
                           gi_5_0_port, P2 => pi_5_0_port, gout => n_1049, pout
                           => n_1050);
   pg_port2_1_7 : PG_38 port map( G1 => gi_7_0_port, P1 => pi_7_0_port, G2 => 
                           gi_6_0_port, P2 => pi_6_0_port, gout => n_1051, pout
                           => n_1052);
   pg_port2_1_8 : PG_37 port map( G1 => gi_8_0_port, P1 => pi_8_0_port, G2 => 
                           gi_7_0_port, P2 => pi_7_0_port, gout => gi_8_1_port,
                           pout => pi_8_1_port);
   pg_port2_1_9 : PG_36 port map( G1 => gi_9_0_port, P1 => pi_9_0_port, G2 => 
                           gi_8_0_port, P2 => pi_8_0_port, gout => n_1053, pout
                           => n_1054);
   pg_port2_1_10 : PG_35 port map( G1 => gi_10_0_port, P1 => pi_10_0_port, G2 
                           => gi_9_0_port, P2 => pi_9_0_port, gout => n_1055, 
                           pout => n_1056);
   pg_port2_1_11 : PG_34 port map( G1 => gi_11_0_port, P1 => pi_11_0_port, G2 
                           => gi_10_0_port, P2 => pi_10_0_port, gout => n_1057,
                           pout => n_1058);
   pg_port2_1_12 : PG_33 port map( G1 => gi_12_0_port, P1 => pi_12_0_port, G2 
                           => gi_11_0_port, P2 => pi_11_0_port, gout => 
                           gi_12_1_port, pout => pi_12_1_port);
   pg_port2_1_13 : PG_32 port map( G1 => gi_13_0_port, P1 => pi_13_0_port, G2 
                           => gi_12_0_port, P2 => pi_12_0_port, gout => n_1059,
                           pout => n_1060);
   pg_port2_1_14 : PG_31 port map( G1 => gi_14_0_port, P1 => pi_14_0_port, G2 
                           => gi_13_0_port, P2 => pi_13_0_port, gout => n_1061,
                           pout => n_1062);
   pg_port2_1_15 : PG_30 port map( G1 => gi_15_0_port, P1 => pi_15_0_port, G2 
                           => gi_14_0_port, P2 => pi_14_0_port, gout => n_1063,
                           pout => n_1064);
   pg_port2_1_16 : PG_29 port map( G1 => gi_16_0_port, P1 => pi_16_0_port, G2 
                           => gi_15_0_port, P2 => pi_15_0_port, gout => 
                           gi_16_1_port, pout => pi_16_1_port);
   pg_port2_1_17 : PG_28 port map( G1 => gi_17_0_port, P1 => pi_17_0_port, G2 
                           => gi_16_0_port, P2 => pi_16_0_port, gout => n_1065,
                           pout => n_1066);
   pg_port2_1_18 : PG_27 port map( G1 => gi_18_0_port, P1 => pi_18_0_port, G2 
                           => gi_17_0_port, P2 => pi_17_0_port, gout => n_1067,
                           pout => n_1068);
   pg_port2_1_19 : PG_26 port map( G1 => gi_19_0_port, P1 => pi_19_0_port, G2 
                           => gi_18_0_port, P2 => pi_18_0_port, gout => n_1069,
                           pout => n_1070);
   pg_port2_1_20 : PG_25 port map( G1 => gi_20_0_port, P1 => pi_20_0_port, G2 
                           => gi_19_0_port, P2 => pi_19_0_port, gout => 
                           gi_20_1_port, pout => pi_20_1_port);
   pg_port2_1_21 : PG_24 port map( G1 => gi_21_0_port, P1 => pi_21_0_port, G2 
                           => gi_20_0_port, P2 => pi_20_0_port, gout => n_1071,
                           pout => n_1072);
   pg_port2_1_22 : PG_23 port map( G1 => gi_22_0_port, P1 => pi_22_0_port, G2 
                           => gi_21_0_port, P2 => pi_21_0_port, gout => n_1073,
                           pout => n_1074);
   pg_port2_1_23 : PG_22 port map( G1 => gi_23_0_port, P1 => pi_23_0_port, G2 
                           => gi_22_0_port, P2 => pi_22_0_port, gout => n_1075,
                           pout => n_1076);
   pg_port2_1_24 : PG_21 port map( G1 => gi_24_0_port, P1 => pi_24_0_port, G2 
                           => gi_23_0_port, P2 => pi_23_0_port, gout => 
                           gi_24_1_port, pout => pi_24_1_port);
   pg_port2_1_25 : PG_20 port map( G1 => gi_25_0_port, P1 => pi_25_0_port, G2 
                           => gi_24_0_port, P2 => pi_24_0_port, gout => n_1077,
                           pout => n_1078);
   pg_port2_1_26 : PG_19 port map( G1 => gi_26_0_port, P1 => pi_26_0_port, G2 
                           => gi_25_0_port, P2 => pi_25_0_port, gout => n_1079,
                           pout => n_1080);
   pg_port2_1_27 : PG_18 port map( G1 => gi_27_0_port, P1 => pi_27_0_port, G2 
                           => gi_26_0_port, P2 => pi_26_0_port, gout => n_1081,
                           pout => n_1082);
   pg_port2_1_28 : PG_17 port map( G1 => gi_28_0_port, P1 => pi_28_0_port, G2 
                           => gi_27_0_port, P2 => pi_27_0_port, gout => 
                           gi_28_1_port, pout => pi_28_1_port);
   pg_port2_1_29 : PG_16 port map( G1 => gi_29_0_port, P1 => pi_29_0_port, G2 
                           => gi_28_0_port, P2 => pi_28_0_port, gout => n_1083,
                           pout => n_1084);
   pg_port2_1_30 : PG_15 port map( G1 => gi_30_0_port, P1 => pi_30_0_port, G2 
                           => gi_29_0_port, P2 => pi_29_0_port, gout => n_1085,
                           pout => n_1086);
   pg_port2_1_31 : PG_14 port map( G1 => gi_31_0_port, P1 => pi_31_0_port, G2 
                           => gi_30_0_port, P2 => pi_30_0_port, gout => n_1087,
                           pout => n_1088);
   pg_port2_1_32 : PG_13 port map( G1 => gi_32_0_port, P1 => pi_32_0_port, G2 
                           => gi_31_0_port, P2 => pi_31_0_port, gout => 
                           gi_32_1_port, pout => pi_32_1_port);
   g_port_0 : G_51 port map( G1 => gi_4_1_port, P => pi_4_1_port, G2 => 
                           gi_2_1_port, Co => Co_0_port);
   pg_port2_0_1_2 : PG_12 port map( G1 => gi_8_1_port, P1 => pi_8_1_port, G2 =>
                           gi_4_1_port, P2 => pi_4_1_port, gout => gi_8_2_port,
                           pout => pi_8_2_port);
   pg_port2_0_2_3 : PG_11 port map( G1 => gi_12_1_port, P1 => pi_12_1_port, G2 
                           => gi_8_1_port, P2 => pi_8_1_port, gout => 
                           gi_12_2_port, pout => pi_12_2_port);
   pg_port2_0_3_4 : PG_10 port map( G1 => gi_16_1_port, P1 => pi_16_1_port, G2 
                           => gi_12_1_port, P2 => pi_12_1_port, gout => 
                           gi_16_2_port, pout => pi_16_2_port);
   pg_port2_0_4_5 : PG_9 port map( G1 => gi_20_1_port, P1 => pi_20_1_port, G2 
                           => gi_16_1_port, P2 => pi_16_1_port, gout => 
                           gi_20_2_port, pout => pi_20_2_port);
   pg_port2_0_5_6 : PG_8 port map( G1 => gi_24_1_port, P1 => pi_24_1_port, G2 
                           => gi_20_1_port, P2 => pi_20_1_port, gout => 
                           gi_24_2_port, pout => pi_24_2_port);
   pg_port2_0_6_7 : PG_7 port map( G1 => gi_28_1_port, P1 => pi_28_1_port, G2 
                           => gi_24_1_port, P2 => pi_24_1_port, gout => 
                           gi_28_2_port, pout => pi_28_2_port);
   pg_port2_0_7_8 : PG_6 port map( G1 => gi_32_1_port, P1 => pi_32_1_port, G2 
                           => gi_28_1_port, P2 => pi_28_1_port, gout => 
                           gi_32_2_port, pout => pi_32_2_port);
   g_port_1_2 : G_50 port map( G1 => gi_8_2_port, P => pi_8_2_port, G2 => 
                           Co_0_port, Co => Co_1_port);
   pg_port2_1_1_4 : PG_5 port map( G1 => gi_16_2_port, P1 => pi_16_2_port, G2 
                           => gi_12_2_port, P2 => pi_12_2_port, gout => 
                           gi_16_3_port, pout => pi_16_3_port);
   pg_port2_1_2_6 : PG_4 port map( G1 => gi_24_2_port, P1 => pi_24_2_port, G2 
                           => gi_20_2_port, P2 => pi_20_2_port, gout => 
                           gi_24_3_port, pout => pi_24_3_port);
   pg_port2_1_3_8 : PG_3 port map( G1 => gi_32_2_port, P1 => pi_32_2_port, G2 
                           => gi_28_2_port, P2 => pi_28_2_port, gout => 
                           gi_32_3_port, pout => pi_32_3_port);
   g_port_2_3 : G_49 port map( G1 => gi_12_2_port, P => pi_12_2_port, G2 => 
                           Co_1_port, Co => Co_2_port);
   g_port_2_4 : G_48 port map( G1 => gi_16_3_port, P => pi_16_3_port, G2 => 
                           Co_1_port, Co => Co_3_port);
   pg_port2_2_1_7 : PG_2 port map( G1 => gi_28_2_port, P1 => pi_28_2_port, G2 
                           => gi_24_3_port, P2 => pi_24_3_port, gout => 
                           gi_28_4_port, pout => pi_28_4_port);
   pg_port2_2_1_8 : PG_1 port map( G1 => gi_32_3_port, P1 => pi_32_3_port, G2 
                           => gi_24_3_port, P2 => pi_24_3_port, gout => 
                           gi_32_4_port, pout => pi_32_4_port);
   g_port_3_5 : G_47 port map( G1 => gi_20_2_port, P => pi_20_2_port, G2 => 
                           Co_3_port, Co => Co_4_port);
   g_port_3_6 : G_46 port map( G1 => gi_24_3_port, P => pi_24_3_port, G2 => 
                           Co_3_port, Co => Co_5_port);
   g_port_3_7 : G_45 port map( G1 => gi_28_4_port, P => pi_28_4_port, G2 => 
                           Co_3_port, Co => Co_6_port);
   g_port_3_8 : G_44 port map( G1 => gi_32_4_port, P => pi_32_4_port, G2 => 
                           Co_3_port, Co => Co_7_port);
   U2 : AND2_X1 port map( A1 => B(31), A2 => A(31), ZN => gi_32_0_port);
   U3 : AND2_X1 port map( A1 => B(15), A2 => A(15), ZN => gi_16_0_port);
   U4 : AND2_X1 port map( A1 => B(14), A2 => A(14), ZN => gi_15_0_port);
   U5 : AND2_X1 port map( A1 => B(19), A2 => A(19), ZN => gi_20_0_port);
   U6 : AND2_X1 port map( A1 => B(18), A2 => A(18), ZN => gi_19_0_port);
   U7 : AND2_X1 port map( A1 => B(23), A2 => A(23), ZN => gi_24_0_port);
   U8 : AND2_X1 port map( A1 => B(22), A2 => A(22), ZN => gi_23_0_port);
   U9 : AND2_X1 port map( A1 => B(27), A2 => A(27), ZN => gi_28_0_port);
   U10 : AND2_X1 port map( A1 => B(26), A2 => A(26), ZN => gi_27_0_port);
   U11 : AND2_X1 port map( A1 => B(30), A2 => A(30), ZN => gi_31_0_port);
   U12 : AND2_X1 port map( A1 => B(7), A2 => A(7), ZN => gi_8_0_port);
   U13 : AND2_X1 port map( A1 => B(6), A2 => A(6), ZN => gi_7_0_port);
   U14 : AND2_X1 port map( A1 => B(11), A2 => A(11), ZN => gi_12_0_port);
   U15 : AND2_X1 port map( A1 => B(10), A2 => A(10), ZN => gi_11_0_port);
   U16 : AND2_X1 port map( A1 => B(3), A2 => A(3), ZN => gi_4_0_port);
   U17 : AND2_X1 port map( A1 => B(2), A2 => A(2), ZN => gi_3_0_port);
   U18 : AND2_X1 port map( A1 => B(0), A2 => A(0), ZN => gi_0_0_port);
   U19 : AND2_X1 port map( A1 => B(1), A2 => A(1), ZN => gi_2_0_port);
   U20 : AND2_X1 port map( A1 => B(4), A2 => A(4), ZN => gi_5_0_port);
   U21 : AND2_X1 port map( A1 => B(5), A2 => A(5), ZN => gi_6_0_port);
   U22 : AND2_X1 port map( A1 => B(8), A2 => A(8), ZN => gi_9_0_port);
   U23 : AND2_X1 port map( A1 => B(9), A2 => A(9), ZN => gi_10_0_port);
   U24 : AND2_X1 port map( A1 => B(12), A2 => A(12), ZN => gi_13_0_port);
   U25 : AND2_X1 port map( A1 => B(13), A2 => A(13), ZN => gi_14_0_port);
   U26 : AND2_X1 port map( A1 => B(16), A2 => A(16), ZN => gi_17_0_port);
   U27 : AND2_X1 port map( A1 => B(17), A2 => A(17), ZN => gi_18_0_port);
   U28 : AND2_X1 port map( A1 => B(20), A2 => A(20), ZN => gi_21_0_port);
   U29 : AND2_X1 port map( A1 => B(21), A2 => A(21), ZN => gi_22_0_port);
   U30 : AND2_X1 port map( A1 => B(24), A2 => A(24), ZN => gi_25_0_port);
   U31 : AND2_X1 port map( A1 => B(25), A2 => A(25), ZN => gi_26_0_port);
   U32 : AND2_X1 port map( A1 => B(28), A2 => A(28), ZN => gi_29_0_port);
   U33 : AND2_X1 port map( A1 => B(29), A2 => A(29), ZN => gi_30_0_port);

end SYN_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ND2_0 is

   port( A, B : in std_logic;  Y : out std_logic);

end ND2_0;

architecture SYN_ARCH2 of ND2_0 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => Y);

end SYN_ARCH2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IV_0 is

   port( A : in std_logic;  Y : out std_logic);

end IV_0;

architecture SYN_BEHAVIORAL of IV_0 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A, ZN => Y);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity P4_ADDER_NBIT32 is

   port( A, B : in std_logic_vector (31 downto 0);  Cin : in std_logic;  S : 
         out std_logic_vector (31 downto 0);  Cout : out std_logic);

end P4_ADDER_NBIT32;

architecture SYN_STRUCTURAL of P4_ADDER_NBIT32 is

   component SUM_GENERATOR_NBIT_PER_BLOCK4_NBLOCKS8
      port( A, B : in std_logic_vector (31 downto 0);  Ci : in std_logic_vector
            (7 downto 0);  S : out std_logic_vector (31 downto 0));
   end component;
   
   component CARRY_GENERATOR_NBIT32_NBIT_PER_BLOCK4
      port( A, B : in std_logic_vector (31 downto 0);  Cin : in std_logic;  Co 
            : out std_logic_vector (7 downto 0));
   end component;
   
   signal Cout_gen_6_port, Cout_gen_5_port, Cout_gen_4_port, Cout_gen_3_port, 
      Cout_gen_2_port, Cout_gen_1_port, Cout_gen_0_port : std_logic;

begin
   
   carry_logic : CARRY_GENERATOR_NBIT32_NBIT_PER_BLOCK4 port map( A(31) => 
                           A(31), A(30) => A(30), A(29) => A(29), A(28) => 
                           A(28), A(27) => A(27), A(26) => A(26), A(25) => 
                           A(25), A(24) => A(24), A(23) => A(23), A(22) => 
                           A(22), A(21) => A(21), A(20) => A(20), A(19) => 
                           A(19), A(18) => A(18), A(17) => A(17), A(16) => 
                           A(16), A(15) => A(15), A(14) => A(14), A(13) => 
                           A(13), A(12) => A(12), A(11) => A(11), A(10) => 
                           A(10), A(9) => A(9), A(8) => A(8), A(7) => A(7), 
                           A(6) => A(6), A(5) => A(5), A(4) => A(4), A(3) => 
                           A(3), A(2) => A(2), A(1) => A(1), A(0) => A(0), 
                           B(31) => B(31), B(30) => B(30), B(29) => B(29), 
                           B(28) => B(28), B(27) => B(27), B(26) => B(26), 
                           B(25) => B(25), B(24) => B(24), B(23) => B(23), 
                           B(22) => B(22), B(21) => B(21), B(20) => B(20), 
                           B(19) => B(19), B(18) => B(18), B(17) => B(17), 
                           B(16) => B(16), B(15) => B(15), B(14) => B(14), 
                           B(13) => B(13), B(12) => B(12), B(11) => B(11), 
                           B(10) => B(10), B(9) => B(9), B(8) => B(8), B(7) => 
                           B(7), B(6) => B(6), B(5) => B(5), B(4) => B(4), B(3)
                           => B(3), B(2) => B(2), B(1) => B(1), B(0) => B(0), 
                           Cin => Cin, Co(7) => Cout, Co(6) => Cout_gen_6_port,
                           Co(5) => Cout_gen_5_port, Co(4) => Cout_gen_4_port, 
                           Co(3) => Cout_gen_3_port, Co(2) => Cout_gen_2_port, 
                           Co(1) => Cout_gen_1_port, Co(0) => Cout_gen_0_port);
   sum_logic : SUM_GENERATOR_NBIT_PER_BLOCK4_NBLOCKS8 port map( A(31) => A(31),
                           A(30) => A(30), A(29) => A(29), A(28) => A(28), 
                           A(27) => A(27), A(26) => A(26), A(25) => A(25), 
                           A(24) => A(24), A(23) => A(23), A(22) => A(22), 
                           A(21) => A(21), A(20) => A(20), A(19) => A(19), 
                           A(18) => A(18), A(17) => A(17), A(16) => A(16), 
                           A(15) => A(15), A(14) => A(14), A(13) => A(13), 
                           A(12) => A(12), A(11) => A(11), A(10) => A(10), A(9)
                           => A(9), A(8) => A(8), A(7) => A(7), A(6) => A(6), 
                           A(5) => A(5), A(4) => A(4), A(3) => A(3), A(2) => 
                           A(2), A(1) => A(1), A(0) => A(0), B(31) => B(31), 
                           B(30) => B(30), B(29) => B(29), B(28) => B(28), 
                           B(27) => B(27), B(26) => B(26), B(25) => B(25), 
                           B(24) => B(24), B(23) => B(23), B(22) => B(22), 
                           B(21) => B(21), B(20) => B(20), B(19) => B(19), 
                           B(18) => B(18), B(17) => B(17), B(16) => B(16), 
                           B(15) => B(15), B(14) => B(14), B(13) => B(13), 
                           B(12) => B(12), B(11) => B(11), B(10) => B(10), B(9)
                           => B(9), B(8) => B(8), B(7) => B(7), B(6) => B(6), 
                           B(5) => B(5), B(4) => B(4), B(3) => B(3), B(2) => 
                           B(2), B(1) => B(1), B(0) => B(0), Ci(7) => 
                           Cout_gen_6_port, Ci(6) => Cout_gen_5_port, Ci(5) => 
                           Cout_gen_4_port, Ci(4) => Cout_gen_3_port, Ci(3) => 
                           Cout_gen_2_port, Ci(2) => Cout_gen_1_port, Ci(1) => 
                           Cout_gen_0_port, Ci(0) => Cin, S(31) => S(31), S(30)
                           => S(30), S(29) => S(29), S(28) => S(28), S(27) => 
                           S(27), S(26) => S(26), S(25) => S(25), S(24) => 
                           S(24), S(23) => S(23), S(22) => S(22), S(21) => 
                           S(21), S(20) => S(20), S(19) => S(19), S(18) => 
                           S(18), S(17) => S(17), S(16) => S(16), S(15) => 
                           S(15), S(14) => S(14), S(13) => S(13), S(12) => 
                           S(12), S(11) => S(11), S(10) => S(10), S(9) => S(9),
                           S(8) => S(8), S(7) => S(7), S(6) => S(6), S(5) => 
                           S(5), S(4) => S(4), S(3) => S(3), S(2) => S(2), S(1)
                           => S(1), S(0) => S(0));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity SHIFTER_GENERIC_N32 is

   port( A : in std_logic_vector (31 downto 0);  B : in std_logic_vector (4 
         downto 0);  LOGIC_ARITH, LEFT_RIGHT, SHIFT_ROTATE : in std_logic;  
         OUTPUT : out std_logic_vector (31 downto 0));

end SHIFTER_GENERIC_N32;

architecture SYN_BEHAVIORAL of SHIFTER_GENERIC_N32 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component SHIFTER_GENERIC_N32_DW_rbsh_0
      port( A : in std_logic_vector (31 downto 0);  SH : in std_logic_vector (4
            downto 0);  SH_TC : in std_logic;  B : out std_logic_vector (31 
            downto 0));
   end component;
   
   component SHIFTER_GENERIC_N32_DW_lbsh_0
      port( A : in std_logic_vector (31 downto 0);  SH : in std_logic_vector (4
            downto 0);  SH_TC : in std_logic;  B : out std_logic_vector (31 
            downto 0));
   end component;
   
   component SHIFTER_GENERIC_N32_DW_sra_0
      port( A : in std_logic_vector (31 downto 0);  SH : in std_logic_vector (4
            downto 0);  SH_TC : in std_logic;  B : out std_logic_vector (31 
            downto 0));
   end component;
   
   component SHIFTER_GENERIC_N32_DW_rash_0
      port( A : in std_logic_vector (31 downto 0);  DATA_TC : in std_logic;  SH
            : in std_logic_vector (4 downto 0);  SH_TC : in std_logic;  B : out
            std_logic_vector (31 downto 0));
   end component;
   
   component SHIFTER_GENERIC_N32_DW_sla_0
      port( A : in std_logic_vector (31 downto 0);  SH : in std_logic_vector (4
            downto 0);  SH_TC : in std_logic;  B : out std_logic_vector (31 
            downto 0));
   end component;
   
   component SHIFTER_GENERIC_N32_DW01_ash_0
      port( A : in std_logic_vector (31 downto 0);  DATA_TC : in std_logic;  SH
            : in std_logic_vector (4 downto 0);  SH_TC : in std_logic;  B : out
            std_logic_vector (31 downto 0));
   end component;
   
   signal N7, N8, N9, N10, N11, N12, N13, N14, N15, N16, N17, N18, N19, N20, 
      N21, N22, N23, N24, N25, N26, N27, N28, N29, N30, N31, N32, N33, N34, N35
      , N36, N37, N38, N39, N40, N41, N42, N43, N44, N45, N46, N47, N48, N49, 
      N50, N51, N52, N53, N54, N55, N56, N57, N58, N59, N60, N61, N62, N63, N64
      , N65, N66, N67, N68, N69, N70, N105, N106, N107, N108, N109, N110, N111,
      N112, N113, N114, N115, N116, N117, N118, N119, N120, N121, N122, N123, 
      N124, N125, N126, N127, N128, N129, N130, N131, N132, N133, N134, N135, 
      N136, N137, N138, N139, N140, N141, N142, N143, N144, N145, N146, N147, 
      N148, N149, N150, N151, N152, N153, N154, N155, N156, N157, N158, N159, 
      N160, N161, N162, N163, N164, N165, N166, N167, N168, N202, N203, N204, 
      N205, N206, N207, N208, N209, N210, N211, N212, N213, N214, N215, N216, 
      N217, N218, N219, N220, N221, N222, N223, N224, N225, N226, N227, N228, 
      N229, N230, N231, N232, N233, N234, N235, N236, N237, N238, N239, N240, 
      N241, N242, N243, N244, N245, N246, N247, N248, N249, N250, N251, N252, 
      N253, N254, N255, N256, N257, N258, N259, N260, N261, N262, N263, N264, 
      N265, n13_port, n14_port, n15_port, n16_port, n17_port, n18_port, 
      n21_port, n22_port, n23_port, n24_port, n25_port, n26_port, n27_port, 
      n28_port, n29_port, n30_port, n31_port, n32_port, n33_port, n34_port, 
      n35_port, n36_port, n37_port, n38_port, n39_port, n40_port, n41_port, 
      n42_port, n43_port, n44_port, n45_port, n46_port, n47_port, n48_port, 
      n49_port, n50_port, n51_port, n52_port, n53_port, n54_port, n55_port, 
      n56_port, n57_port, n58_port, n59_port, n60_port, n61_port, n62_port, 
      n63_port, n64_port, n65_port, n66_port, n67_port, n68_port, n69_port, 
      n70_port, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83
      , n84, n85, n86, n87, n88, n89, n90, n91, n92, n1, n2, n3, n4, n5, n6, 
      n7_port, n8_port, n9_port, n10_port, n11_port, n12_port, n19_port, 
      n20_port, n93, n94, n95, n96, n97, n98, n99 : std_logic;

begin
   
   n13_port <= '0';
   n14_port <= '0';
   n15_port <= '0';
   n16_port <= '0';
   n17_port <= '0';
   n18_port <= '0';
   sll_49 : SHIFTER_GENERIC_N32_DW01_ash_0 port map( A(31) => A(31), A(30) => 
                           A(30), A(29) => A(29), A(28) => A(28), A(27) => 
                           A(27), A(26) => A(26), A(25) => A(25), A(24) => 
                           A(24), A(23) => A(23), A(22) => A(22), A(21) => 
                           A(21), A(20) => A(20), A(19) => A(19), A(18) => 
                           A(18), A(17) => A(17), A(16) => A(16), A(15) => 
                           A(15), A(14) => A(14), A(13) => A(13), A(12) => 
                           A(12), A(11) => A(11), A(10) => A(10), A(9) => A(9),
                           A(8) => A(8), A(7) => A(7), A(6) => A(6), A(5) => 
                           A(5), A(4) => A(4), A(3) => A(3), A(2) => A(2), A(1)
                           => A(1), A(0) => A(0), DATA_TC => n13_port, SH(4) =>
                           n97, SH(3) => B(3), SH(2) => B(2), SH(1) => B(1), 
                           SH(0) => B(0), SH_TC => n13_port, B(31) => N265, 
                           B(30) => N264, B(29) => N263, B(28) => N262, B(27) 
                           => N261, B(26) => N260, B(25) => N259, B(24) => N258
                           , B(23) => N257, B(22) => N256, B(21) => N255, B(20)
                           => N254, B(19) => N253, B(18) => N252, B(17) => N251
                           , B(16) => N250, B(15) => N249, B(14) => N248, B(13)
                           => N247, B(12) => N246, B(11) => N245, B(10) => N244
                           , B(9) => N243, B(8) => N242, B(7) => N241, B(6) => 
                           N240, B(5) => N239, B(4) => N238, B(3) => N237, B(2)
                           => N236, B(1) => N235, B(0) => N234);
   sla_47 : SHIFTER_GENERIC_N32_DW_sla_0 port map( A(31) => A(31), A(30) => 
                           A(30), A(29) => A(29), A(28) => A(28), A(27) => 
                           A(27), A(26) => A(26), A(25) => A(25), A(24) => 
                           A(24), A(23) => A(23), A(22) => A(22), A(21) => 
                           A(21), A(20) => A(20), A(19) => A(19), A(18) => 
                           A(18), A(17) => A(17), A(16) => A(16), A(15) => 
                           A(15), A(14) => A(14), A(13) => A(13), A(12) => 
                           A(12), A(11) => A(11), A(10) => A(10), A(9) => A(9),
                           A(8) => A(8), A(7) => A(7), A(6) => A(6), A(5) => 
                           A(5), A(4) => A(4), A(3) => A(3), A(2) => A(2), A(1)
                           => A(1), A(0) => A(0), SH(4) => n97, SH(3) => B(3), 
                           SH(2) => B(2), SH(1) => B(1), SH(0) => B(0), SH_TC 
                           => n14_port, B(31) => N233, B(30) => N232, B(29) => 
                           N231, B(28) => N230, B(27) => N229, B(26) => N228, 
                           B(25) => N227, B(24) => N226, B(23) => N225, B(22) 
                           => N224, B(21) => N223, B(20) => N222, B(19) => N221
                           , B(18) => N220, B(17) => N219, B(16) => N218, B(15)
                           => N217, B(14) => N216, B(13) => N215, B(12) => N214
                           , B(11) => N213, B(10) => N212, B(9) => N211, B(8) 
                           => N210, B(7) => N209, B(6) => N208, B(5) => N207, 
                           B(4) => N206, B(3) => N205, B(2) => N204, B(1) => 
                           N203, B(0) => N202);
   srl_42 : SHIFTER_GENERIC_N32_DW_rash_0 port map( A(31) => A(31), A(30) => 
                           A(30), A(29) => A(29), A(28) => A(28), A(27) => 
                           A(27), A(26) => A(26), A(25) => A(25), A(24) => 
                           A(24), A(23) => A(23), A(22) => A(22), A(21) => 
                           A(21), A(20) => A(20), A(19) => A(19), A(18) => 
                           A(18), A(17) => A(17), A(16) => A(16), A(15) => 
                           A(15), A(14) => A(14), A(13) => A(13), A(12) => 
                           A(12), A(11) => A(11), A(10) => A(10), A(9) => A(9),
                           A(8) => A(8), A(7) => A(7), A(6) => A(6), A(5) => 
                           A(5), A(4) => A(4), A(3) => A(3), A(2) => A(2), A(1)
                           => A(1), A(0) => A(0), DATA_TC => n15_port, SH(4) =>
                           n97, SH(3) => B(3), SH(2) => B(2), SH(1) => B(1), 
                           SH(0) => B(0), SH_TC => n15_port, B(31) => N168, 
                           B(30) => N167, B(29) => N166, B(28) => N165, B(27) 
                           => N164, B(26) => N163, B(25) => N162, B(24) => N161
                           , B(23) => N160, B(22) => N159, B(21) => N158, B(20)
                           => N157, B(19) => N156, B(18) => N155, B(17) => N154
                           , B(16) => N153, B(15) => N152, B(14) => N151, B(13)
                           => N150, B(12) => N149, B(11) => N148, B(10) => N147
                           , B(9) => N146, B(8) => N145, B(7) => N144, B(6) => 
                           N143, B(5) => N142, B(4) => N141, B(3) => N140, B(2)
                           => N139, B(1) => N138, B(0) => N137);
   sra_40 : SHIFTER_GENERIC_N32_DW_sra_0 port map( A(31) => A(31), A(30) => 
                           A(30), A(29) => A(29), A(28) => A(28), A(27) => 
                           A(27), A(26) => A(26), A(25) => A(25), A(24) => 
                           A(24), A(23) => A(23), A(22) => A(22), A(21) => 
                           A(21), A(20) => A(20), A(19) => A(19), A(18) => 
                           A(18), A(17) => A(17), A(16) => A(16), A(15) => 
                           A(15), A(14) => A(14), A(13) => A(13), A(12) => 
                           A(12), A(11) => A(11), A(10) => A(10), A(9) => A(9),
                           A(8) => A(8), A(7) => A(7), A(6) => A(6), A(5) => 
                           A(5), A(4) => A(4), A(3) => A(3), A(2) => A(2), A(1)
                           => A(1), A(0) => A(0), SH(4) => n97, SH(3) => B(3), 
                           SH(2) => B(2), SH(1) => B(1), SH(0) => B(0), SH_TC 
                           => n16_port, B(31) => N136, B(30) => N135, B(29) => 
                           N134, B(28) => N133, B(27) => N132, B(26) => N131, 
                           B(25) => N130, B(24) => N129, B(23) => N128, B(22) 
                           => N127, B(21) => N126, B(20) => N125, B(19) => N124
                           , B(18) => N123, B(17) => N122, B(16) => N121, B(15)
                           => N120, B(14) => N119, B(13) => N118, B(12) => N117
                           , B(11) => N116, B(10) => N115, B(9) => N114, B(8) 
                           => N113, B(7) => N112, B(6) => N111, B(5) => N110, 
                           B(4) => N109, B(3) => N108, B(2) => N107, B(1) => 
                           N106, B(0) => N105);
   rol_33 : SHIFTER_GENERIC_N32_DW_lbsh_0 port map( A(31) => A(31), A(30) => 
                           A(30), A(29) => A(29), A(28) => A(28), A(27) => 
                           A(27), A(26) => A(26), A(25) => A(25), A(24) => 
                           A(24), A(23) => A(23), A(22) => A(22), A(21) => 
                           A(21), A(20) => A(20), A(19) => A(19), A(18) => 
                           A(18), A(17) => A(17), A(16) => A(16), A(15) => 
                           A(15), A(14) => A(14), A(13) => A(13), A(12) => 
                           A(12), A(11) => A(11), A(10) => A(10), A(9) => A(9),
                           A(8) => A(8), A(7) => A(7), A(6) => A(6), A(5) => 
                           A(5), A(4) => A(4), A(3) => A(3), A(2) => A(2), A(1)
                           => A(1), A(0) => A(0), SH(4) => n97, SH(3) => B(3), 
                           SH(2) => B(2), SH(1) => B(1), SH(0) => B(0), SH_TC 
                           => n17_port, B(31) => N70, B(30) => N69, B(29) => 
                           N68, B(28) => N67, B(27) => N66, B(26) => N65, B(25)
                           => N64, B(24) => N63, B(23) => N62, B(22) => N61, 
                           B(21) => N60, B(20) => N59, B(19) => N58, B(18) => 
                           N57, B(17) => N56, B(16) => N55, B(15) => N54, B(14)
                           => N53, B(13) => N52, B(12) => N51, B(11) => N50, 
                           B(10) => N49, B(9) => N48, B(8) => N47, B(7) => N46,
                           B(6) => N45, B(5) => N44, B(4) => N43, B(3) => N42, 
                           B(2) => N41, B(1) => N40, B(0) => N39);
   ror_31 : SHIFTER_GENERIC_N32_DW_rbsh_0 port map( A(31) => A(31), A(30) => 
                           A(30), A(29) => A(29), A(28) => A(28), A(27) => 
                           A(27), A(26) => A(26), A(25) => A(25), A(24) => 
                           A(24), A(23) => A(23), A(22) => A(22), A(21) => 
                           A(21), A(20) => A(20), A(19) => A(19), A(18) => 
                           A(18), A(17) => A(17), A(16) => A(16), A(15) => 
                           A(15), A(14) => A(14), A(13) => A(13), A(12) => 
                           A(12), A(11) => A(11), A(10) => A(10), A(9) => A(9),
                           A(8) => A(8), A(7) => A(7), A(6) => A(6), A(5) => 
                           A(5), A(4) => A(4), A(3) => A(3), A(2) => A(2), A(1)
                           => A(1), A(0) => A(0), SH(4) => n97, SH(3) => B(3), 
                           SH(2) => B(2), SH(1) => B(1), SH(0) => B(0), SH_TC 
                           => n18_port, B(31) => N38, B(30) => N37, B(29) => 
                           N36, B(28) => N35, B(27) => N34, B(26) => N33, B(25)
                           => N32, B(24) => N31, B(23) => N30, B(22) => N29, 
                           B(21) => N28, B(20) => N27, B(19) => N26, B(18) => 
                           N25, B(17) => N24, B(16) => N23, B(15) => N22, B(14)
                           => N21, B(13) => N20, B(12) => N19, B(11) => N18, 
                           B(10) => N17, B(9) => N16, B(8) => N15, B(7) => N14,
                           B(6) => N13, B(5) => N12, B(4) => N11, B(3) => N10, 
                           B(2) => N9, B(1) => N8, B(0) => N7);
   U5 : AOI222_X1 port map( A1 => N211, A2 => n96, B1 => N114, B2 => n93, C1 =>
                           N146, C2 => n12_port, ZN => n22_port);
   U6 : AOI222_X1 port map( A1 => N210, A2 => n96, B1 => N113, B2 => n93, C1 =>
                           N145, C2 => n12_port, ZN => n30_port);
   U7 : AOI222_X1 port map( A1 => N209, A2 => n96, B1 => N112, B2 => n93, C1 =>
                           N144, C2 => n12_port, ZN => n32_port);
   U8 : AOI222_X1 port map( A1 => N208, A2 => n96, B1 => N111, B2 => n93, C1 =>
                           N143, C2 => n12_port, ZN => n34_port);
   U9 : AOI222_X1 port map( A1 => N207, A2 => n96, B1 => N110, B2 => n93, C1 =>
                           N142, C2 => n12_port, ZN => n36_port);
   U10 : AOI222_X1 port map( A1 => N206, A2 => n96, B1 => N109, B2 => n93, C1 
                           => N141, C2 => n12_port, ZN => n38_port);
   U13 : AOI222_X1 port map( A1 => N205, A2 => n96, B1 => N108, B2 => n93, C1 
                           => N140, C2 => n12_port, ZN => n40_port);
   U14 : AOI222_X1 port map( A1 => N232, A2 => n95, B1 => N135, B2 => n20_port,
                           C1 => N167, C2 => n11_port, ZN => n44_port);
   U15 : AOI222_X1 port map( A1 => N231, A2 => n95, B1 => N134, B2 => n20_port,
                           C1 => N166, C2 => n11_port, ZN => n48_port);
   U16 : AOI222_X1 port map( A1 => N230, A2 => n95, B1 => N133, B2 => n20_port,
                           C1 => N165, C2 => n11_port, ZN => n50_port);
   U17 : AOI222_X1 port map( A1 => N229, A2 => n95, B1 => N132, B2 => n20_port,
                           C1 => N164, C2 => n11_port, ZN => n52_port);
   U18 : AOI222_X1 port map( A1 => N228, A2 => n95, B1 => N131, B2 => n20_port,
                           C1 => N163, C2 => n11_port, ZN => n54_port);
   U19 : AOI222_X1 port map( A1 => N227, A2 => n95, B1 => N130, B2 => n20_port,
                           C1 => N162, C2 => n11_port, ZN => n56_port);
   U20 : AOI222_X1 port map( A1 => N226, A2 => n95, B1 => N129, B2 => n20_port,
                           C1 => N161, C2 => n11_port, ZN => n58_port);
   U21 : AOI222_X1 port map( A1 => N225, A2 => n95, B1 => N128, B2 => n20_port,
                           C1 => N160, C2 => n11_port, ZN => n60_port);
   U22 : AOI222_X1 port map( A1 => N224, A2 => n95, B1 => N127, B2 => n20_port,
                           C1 => N159, C2 => n11_port, ZN => n62_port);
   U23 : AOI222_X1 port map( A1 => N223, A2 => n95, B1 => N126, B2 => n20_port,
                           C1 => N158, C2 => n11_port, ZN => n64_port);
   U24 : AOI222_X1 port map( A1 => N222, A2 => n95, B1 => N125, B2 => n20_port,
                           C1 => N157, C2 => n11_port, ZN => n66_port);
   U25 : AOI222_X1 port map( A1 => N221, A2 => n94, B1 => N124, B2 => n19_port,
                           C1 => N156, C2 => n10_port, ZN => n70_port);
   U26 : AOI222_X1 port map( A1 => N220, A2 => n94, B1 => N123, B2 => n19_port,
                           C1 => N155, C2 => n10_port, ZN => n72);
   U27 : AOI222_X1 port map( A1 => N219, A2 => n94, B1 => N122, B2 => n19_port,
                           C1 => N154, C2 => n10_port, ZN => n74);
   U28 : AOI222_X1 port map( A1 => N218, A2 => n94, B1 => N121, B2 => n19_port,
                           C1 => N153, C2 => n10_port, ZN => n76);
   U29 : AOI222_X1 port map( A1 => N217, A2 => n94, B1 => N120, B2 => n19_port,
                           C1 => N152, C2 => n10_port, ZN => n78);
   U30 : AOI222_X1 port map( A1 => N216, A2 => n94, B1 => N119, B2 => n19_port,
                           C1 => N151, C2 => n10_port, ZN => n80);
   U31 : AOI222_X1 port map( A1 => N215, A2 => n94, B1 => N118, B2 => n19_port,
                           C1 => N150, C2 => n10_port, ZN => n82);
   U32 : AOI222_X1 port map( A1 => N214, A2 => n94, B1 => N117, B2 => n19_port,
                           C1 => N149, C2 => n10_port, ZN => n84);
   U33 : AOI222_X1 port map( A1 => N213, A2 => n94, B1 => N116, B2 => n19_port,
                           C1 => N148, C2 => n10_port, ZN => n86);
   U34 : AOI222_X1 port map( A1 => N212, A2 => n94, B1 => N115, B2 => n19_port,
                           C1 => N147, C2 => n10_port, ZN => n88);
   U35 : AOI222_X1 port map( A1 => N204, A2 => n95, B1 => N107, B2 => n20_port,
                           C1 => N139, C2 => n11_port, ZN => n46_port);
   U36 : AOI222_X1 port map( A1 => N203, A2 => n94, B1 => N106, B2 => n19_port,
                           C1 => N138, C2 => n10_port, ZN => n68_port);
   U37 : AOI222_X1 port map( A1 => N70, A2 => n9_port, B1 => N265, B2 => n6, C1
                           => N38, C2 => n3, ZN => n41_port);
   U38 : AOI222_X1 port map( A1 => N48, A2 => n9_port, B1 => N243, B2 => n6, C1
                           => N16, C2 => n3, ZN => n21_port);
   U39 : AOI222_X1 port map( A1 => N47, A2 => n9_port, B1 => N242, B2 => n6, C1
                           => N15, C2 => n3, ZN => n29_port);
   U40 : AOI222_X1 port map( A1 => N46, A2 => n9_port, B1 => N241, B2 => n6, C1
                           => N14, C2 => n3, ZN => n31_port);
   U41 : AOI222_X1 port map( A1 => N45, A2 => n9_port, B1 => N240, B2 => n6, C1
                           => N13, C2 => n3, ZN => n33_port);
   U42 : AOI222_X1 port map( A1 => N44, A2 => n9_port, B1 => N239, B2 => n6, C1
                           => N12, C2 => n3, ZN => n35_port);
   U43 : AOI222_X1 port map( A1 => N43, A2 => n9_port, B1 => N238, B2 => n6, C1
                           => N11, C2 => n3, ZN => n37_port);
   U44 : AOI222_X1 port map( A1 => N42, A2 => n9_port, B1 => N237, B2 => n6, C1
                           => N10, C2 => n3, ZN => n39_port);
   U45 : AOI222_X1 port map( A1 => N69, A2 => n8_port, B1 => N264, B2 => n5, C1
                           => N37, C2 => n2, ZN => n43_port);
   U46 : AOI222_X1 port map( A1 => N68, A2 => n8_port, B1 => N263, B2 => n5, C1
                           => N36, C2 => n2, ZN => n47_port);
   U47 : AOI222_X1 port map( A1 => N67, A2 => n8_port, B1 => N262, B2 => n5, C1
                           => N35, C2 => n2, ZN => n49_port);
   U48 : AOI222_X1 port map( A1 => N66, A2 => n8_port, B1 => N261, B2 => n5, C1
                           => N34, C2 => n2, ZN => n51_port);
   U49 : AOI222_X1 port map( A1 => N65, A2 => n8_port, B1 => N260, B2 => n5, C1
                           => N33, C2 => n2, ZN => n53_port);
   U50 : AOI222_X1 port map( A1 => N64, A2 => n8_port, B1 => N259, B2 => n5, C1
                           => N32, C2 => n2, ZN => n55_port);
   U51 : AOI222_X1 port map( A1 => N63, A2 => n8_port, B1 => N258, B2 => n5, C1
                           => N31, C2 => n2, ZN => n57_port);
   U52 : AOI222_X1 port map( A1 => N62, A2 => n8_port, B1 => N257, B2 => n5, C1
                           => N30, C2 => n2, ZN => n59_port);
   U53 : AOI222_X1 port map( A1 => N61, A2 => n8_port, B1 => N256, B2 => n5, C1
                           => N29, C2 => n2, ZN => n61_port);
   U54 : AOI222_X1 port map( A1 => N60, A2 => n8_port, B1 => N255, B2 => n5, C1
                           => N28, C2 => n2, ZN => n63_port);
   U55 : AOI222_X1 port map( A1 => N59, A2 => n8_port, B1 => N254, B2 => n5, C1
                           => N27, C2 => n2, ZN => n65_port);
   U56 : AOI222_X1 port map( A1 => N58, A2 => n7_port, B1 => N253, B2 => n4, C1
                           => N26, C2 => n1, ZN => n69_port);
   U57 : AOI222_X1 port map( A1 => N57, A2 => n7_port, B1 => N252, B2 => n4, C1
                           => N25, C2 => n1, ZN => n71);
   U58 : AOI222_X1 port map( A1 => N56, A2 => n7_port, B1 => N251, B2 => n4, C1
                           => N24, C2 => n1, ZN => n73);
   U59 : AOI222_X1 port map( A1 => N55, A2 => n7_port, B1 => N250, B2 => n4, C1
                           => N23, C2 => n1, ZN => n75);
   U60 : AOI222_X1 port map( A1 => N54, A2 => n7_port, B1 => N249, B2 => n4, C1
                           => N22, C2 => n1, ZN => n77);
   U61 : AOI222_X1 port map( A1 => N53, A2 => n7_port, B1 => N248, B2 => n4, C1
                           => N21, C2 => n1, ZN => n79);
   U62 : AOI222_X1 port map( A1 => N52, A2 => n7_port, B1 => N247, B2 => n4, C1
                           => N20, C2 => n1, ZN => n81);
   U63 : AOI222_X1 port map( A1 => N51, A2 => n7_port, B1 => N246, B2 => n4, C1
                           => N19, C2 => n1, ZN => n83);
   U64 : AOI222_X1 port map( A1 => N50, A2 => n7_port, B1 => N245, B2 => n4, C1
                           => N18, C2 => n1, ZN => n85);
   U65 : AOI222_X1 port map( A1 => N49, A2 => n7_port, B1 => N244, B2 => n4, C1
                           => N17, C2 => n1, ZN => n87);
   U66 : AOI222_X1 port map( A1 => N41, A2 => n8_port, B1 => N236, B2 => n5, C1
                           => N9, C2 => n2, ZN => n45_port);
   U67 : AOI222_X1 port map( A1 => N40, A2 => n7_port, B1 => N235, B2 => n4, C1
                           => N8, C2 => n1, ZN => n67_port);
   U68 : AOI222_X1 port map( A1 => N39, A2 => n7_port, B1 => N234, B2 => n4, C1
                           => N7, C2 => n1, ZN => n89);
   U69 : BUF_X1 port map( A => n24_port, Z => n20_port);
   U70 : BUF_X1 port map( A => n24_port, Z => n19_port);
   U71 : BUF_X1 port map( A => n25_port, Z => n11_port);
   U72 : BUF_X1 port map( A => n25_port, Z => n10_port);
   U73 : BUF_X1 port map( A => n24_port, Z => n93);
   U74 : BUF_X1 port map( A => n25_port, Z => n12_port);
   U75 : BUF_X1 port map( A => B(4), Z => n97);
   U76 : NAND2_X1 port map( A1 => n41_port, A2 => n42_port, ZN => OUTPUT(31));
   U77 : NAND2_X1 port map( A1 => n43_port, A2 => n44_port, ZN => OUTPUT(30));
   U78 : NAND2_X1 port map( A1 => n47_port, A2 => n48_port, ZN => OUTPUT(29));
   U79 : NAND2_X1 port map( A1 => n49_port, A2 => n50_port, ZN => OUTPUT(28));
   U80 : NAND2_X1 port map( A1 => n51_port, A2 => n52_port, ZN => OUTPUT(27));
   U81 : NAND2_X1 port map( A1 => n53_port, A2 => n54_port, ZN => OUTPUT(26));
   U82 : NAND2_X1 port map( A1 => n55_port, A2 => n56_port, ZN => OUTPUT(25));
   U83 : NAND2_X1 port map( A1 => n57_port, A2 => n58_port, ZN => OUTPUT(24));
   U84 : NAND2_X1 port map( A1 => n59_port, A2 => n60_port, ZN => OUTPUT(23));
   U85 : NAND2_X1 port map( A1 => n61_port, A2 => n62_port, ZN => OUTPUT(22));
   U86 : NAND2_X1 port map( A1 => n63_port, A2 => n64_port, ZN => OUTPUT(21));
   U87 : NAND2_X1 port map( A1 => n65_port, A2 => n66_port, ZN => OUTPUT(20));
   U88 : NAND2_X1 port map( A1 => n69_port, A2 => n70_port, ZN => OUTPUT(19));
   U89 : NAND2_X1 port map( A1 => n71, A2 => n72, ZN => OUTPUT(18));
   U90 : NAND2_X1 port map( A1 => n73, A2 => n74, ZN => OUTPUT(17));
   U91 : NAND2_X1 port map( A1 => n75, A2 => n76, ZN => OUTPUT(16));
   U92 : NAND2_X1 port map( A1 => n77, A2 => n78, ZN => OUTPUT(15));
   U93 : NAND2_X1 port map( A1 => n79, A2 => n80, ZN => OUTPUT(14));
   U94 : NAND2_X1 port map( A1 => n81, A2 => n82, ZN => OUTPUT(13));
   U95 : NAND2_X1 port map( A1 => n83, A2 => n84, ZN => OUTPUT(12));
   U96 : NAND2_X1 port map( A1 => n85, A2 => n86, ZN => OUTPUT(11));
   U97 : NAND2_X1 port map( A1 => n87, A2 => n88, ZN => OUTPUT(10));
   U98 : NAND2_X1 port map( A1 => n21_port, A2 => n22_port, ZN => OUTPUT(9));
   U99 : NAND2_X1 port map( A1 => n29_port, A2 => n30_port, ZN => OUTPUT(8));
   U100 : NAND2_X1 port map( A1 => n31_port, A2 => n32_port, ZN => OUTPUT(7));
   U101 : NAND2_X1 port map( A1 => n33_port, A2 => n34_port, ZN => OUTPUT(6));
   U102 : NAND2_X1 port map( A1 => n35_port, A2 => n36_port, ZN => OUTPUT(5));
   U103 : NAND2_X1 port map( A1 => n37_port, A2 => n38_port, ZN => OUTPUT(4));
   U104 : AOI222_X1 port map( A1 => N233, A2 => n96, B1 => N136, B2 => n93, C1 
                           => N168, C2 => n12_port, ZN => n42_port);
   U105 : AOI222_X1 port map( A1 => N202, A2 => n94, B1 => N105, B2 => n19_port
                           , C1 => N137, C2 => n10_port, ZN => n90);
   U106 : BUF_X1 port map( A => n27_port, Z => n5);
   U107 : BUF_X1 port map( A => n27_port, Z => n4);
   U108 : BUF_X1 port map( A => n28_port, Z => n2);
   U109 : BUF_X1 port map( A => n28_port, Z => n1);
   U110 : BUF_X1 port map( A => n26_port, Z => n8_port);
   U111 : BUF_X1 port map( A => n26_port, Z => n7_port);
   U112 : BUF_X1 port map( A => n23_port, Z => n95);
   U113 : BUF_X1 port map( A => n23_port, Z => n94);
   U114 : BUF_X1 port map( A => n27_port, Z => n6);
   U115 : BUF_X1 port map( A => n28_port, Z => n3);
   U116 : BUF_X1 port map( A => n26_port, Z => n9_port);
   U117 : BUF_X1 port map( A => n23_port, Z => n96);
   U118 : AND2_X1 port map( A1 => n92, A2 => n98, ZN => n24_port);
   U119 : AND2_X1 port map( A1 => n91, A2 => n98, ZN => n25_port);
   U120 : NAND2_X1 port map( A1 => n39_port, A2 => n40_port, ZN => OUTPUT(3));
   U121 : NAND2_X1 port map( A1 => n45_port, A2 => n46_port, ZN => OUTPUT(2));
   U122 : NAND2_X1 port map( A1 => n67_port, A2 => n68_port, ZN => OUTPUT(1));
   U123 : NOR2_X1 port map( A1 => LEFT_RIGHT, A2 => SHIFT_ROTATE, ZN => 
                           n28_port);
   U124 : NOR2_X1 port map( A1 => n98, A2 => SHIFT_ROTATE, ZN => n26_port);
   U125 : NOR2_X1 port map( A1 => n99, A2 => LOGIC_ARITH, ZN => n92);
   U126 : INV_X1 port map( A => SHIFT_ROTATE, ZN => n99);
   U127 : AND2_X1 port map( A1 => LEFT_RIGHT, A2 => n92, ZN => n23_port);
   U128 : AND2_X1 port map( A1 => LEFT_RIGHT, A2 => n91, ZN => n27_port);
   U129 : INV_X1 port map( A => LEFT_RIGHT, ZN => n98);
   U130 : AND2_X1 port map( A1 => LOGIC_ARITH, A2 => SHIFT_ROTATE, ZN => n91);
   U131 : NAND2_X1 port map( A1 => n89, A2 => n90, ZN => OUTPUT(0));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity comparator is

   port( DATA1 : in std_logic_vector (31 downto 0);  DATA2i : in std_logic;  
         tipo : in std_logic_vector (0 to 5);  OUTALU : out std_logic_vector 
         (31 downto 0));

end comparator;

architecture SYN_Architectural of comparator is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N57, N58, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23,
      n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38
      , n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n1, n2, n3, n4, 
      n5, n6, n7, n8, n9, n10, n11 : std_logic;

begin
   
   OUTALU_reg_0_inst : DLH_X1 port map( G => N57, D => N58, Q => OUTALU(0));
   OUTALU(1) <= '0';
   OUTALU(2) <= '0';
   OUTALU(3) <= '0';
   OUTALU(4) <= '0';
   OUTALU(5) <= '0';
   OUTALU(6) <= '0';
   OUTALU(7) <= '0';
   OUTALU(8) <= '0';
   OUTALU(9) <= '0';
   OUTALU(10) <= '0';
   OUTALU(11) <= '0';
   OUTALU(12) <= '0';
   OUTALU(13) <= '0';
   OUTALU(14) <= '0';
   OUTALU(15) <= '0';
   OUTALU(16) <= '0';
   OUTALU(17) <= '0';
   OUTALU(18) <= '0';
   OUTALU(19) <= '0';
   OUTALU(20) <= '0';
   OUTALU(21) <= '0';
   OUTALU(22) <= '0';
   OUTALU(23) <= '0';
   OUTALU(24) <= '0';
   OUTALU(25) <= '0';
   OUTALU(26) <= '0';
   OUTALU(27) <= '0';
   OUTALU(28) <= '0';
   OUTALU(29) <= '0';
   OUTALU(30) <= '0';
   OUTALU(31) <= '0';
   U80 : NAND3_X1 port map( A1 => n48, A2 => n7, A3 => tipo(0), ZN => n37);
   U81 : NAND3_X1 port map( A1 => tipo(2), A2 => n48, A3 => tipo(0), ZN => n43)
                           ;
   U82 : NAND3_X1 port map( A1 => tipo(2), A2 => n49, A3 => tipo(4), ZN => n46)
                           ;
   U83 : NAND3_X1 port map( A1 => n48, A2 => n5, A3 => tipo(2), ZN => n42);
   U33 : INV_X1 port map( A => n19, ZN => n1);
   U34 : NOR4_X1 port map( A1 => DATA1(23), A2 => DATA1(22), A3 => DATA1(21), 
                           A4 => DATA1(20), ZN => n27);
   U35 : NOR4_X1 port map( A1 => DATA1(9), A2 => DATA1(8), A3 => DATA1(7), A4 
                           => DATA1(6), ZN => n31);
   U36 : NOR4_X1 port map( A1 => DATA1(16), A2 => DATA1(15), A3 => DATA1(14), 
                           A4 => DATA1(13), ZN => n25);
   U37 : NOR2_X1 port map( A1 => n22, A2 => n23, ZN => n19);
   U38 : NAND4_X1 port map( A1 => n28, A2 => n29, A3 => n30, A4 => n31, ZN => 
                           n22);
   U39 : NAND4_X1 port map( A1 => n24, A2 => n25, A3 => n26, A4 => n27, ZN => 
                           n23);
   U40 : NOR4_X1 port map( A1 => DATA1(27), A2 => DATA1(26), A3 => DATA1(25), 
                           A4 => DATA1(24), ZN => n28);
   U41 : INV_X1 port map( A => DATA2i, ZN => n2);
   U42 : NOR4_X1 port map( A1 => DATA1(1), A2 => DATA1(19), A3 => DATA1(18), A4
                           => DATA1(17), ZN => n26);
   U43 : NOR4_X1 port map( A1 => DATA1(5), A2 => DATA1(4), A3 => DATA1(3), A4 
                           => DATA1(31), ZN => n30);
   U44 : NOR4_X1 port map( A1 => DATA1(30), A2 => DATA1(2), A3 => DATA1(29), A4
                           => DATA1(28), ZN => n29);
   U45 : OAI221_X1 port map( B1 => n39, B2 => n36, C1 => n34, C2 => n40, A => 
                           n4, ZN => n21);
   U46 : INV_X1 port map( A => n41, ZN => n4);
   U47 : AOI211_X1 port map( C1 => n37, C2 => n42, A => n9, B => n11, ZN => n41
                           );
   U48 : NOR4_X1 port map( A1 => DATA1(12), A2 => DATA1(11), A3 => DATA1(10), 
                           A4 => DATA1(0), ZN => n24);
   U49 : OAI22_X1 port map( A1 => n39, A2 => n40, B1 => n34, B2 => n42, ZN => 
                           n18);
   U50 : OAI22_X1 port map( A1 => n42, A2 => n39, B1 => n40, B2 => n38, ZN => 
                           n16);
   U51 : OAI21_X1 port map( B1 => n33, B2 => n34, A => n6, ZN => n20);
   U52 : INV_X1 port map( A => n35, ZN => n6);
   U53 : AOI21_X1 port map( B1 => n36, B2 => n37, A => n38, ZN => n35);
   U54 : NAND2_X1 port map( A1 => n11, A2 => n9, ZN => n38);
   U55 : OAI211_X1 port map( C1 => n12, C2 => n2, A => n13, B => n14, ZN => N58
                           );
   U56 : OAI21_X1 port map( B1 => n17, B2 => n18, A => n19, ZN => n13);
   U57 : AOI21_X1 port map( B1 => n20, B2 => n1, A => n21, ZN => n12);
   U58 : AOI22_X1 port map( A1 => n15, A2 => n2, B1 => n16, B2 => n1, ZN => n14
                           );
   U59 : OR4_X1 port map( A1 => n16, A2 => n15, A3 => n32, A4 => n20, ZN => N57
                           );
   U60 : OR2_X1 port map( A1 => n17, A2 => n21, ZN => n32);
   U61 : AND2_X1 port map( A1 => n43, A2 => n37, ZN => n33);
   U62 : NAND4_X1 port map( A1 => tipo(1), A2 => tipo(3), A3 => n7, A4 => n5, 
                           ZN => n40);
   U63 : OAI221_X1 port map( B1 => n46, B2 => n47, C1 => n33, C2 => n39, A => 
                           n3, ZN => n15);
   U64 : INV_X1 port map( A => n18, ZN => n3);
   U65 : NAND2_X1 port map( A1 => tipo(5), A2 => tipo(3), ZN => n47);
   U66 : NAND4_X1 port map( A1 => tipo(0), A2 => tipo(1), A3 => n8, A4 => n7, 
                           ZN => n36);
   U67 : INV_X1 port map( A => tipo(3), ZN => n8);
   U68 : NAND2_X1 port map( A1 => tipo(4), A2 => n11, ZN => n34);
   U69 : NAND2_X1 port map( A1 => tipo(5), A2 => n9, ZN => n39);
   U70 : INV_X1 port map( A => tipo(2), ZN => n7);
   U71 : NOR2_X1 port map( A1 => tipo(1), A2 => tipo(3), ZN => n48);
   U72 : OAI21_X1 port map( B1 => n43, B2 => n38, A => n44, ZN => n17);
   U73 : NAND4_X1 port map( A1 => tipo(1), A2 => tipo(3), A3 => n45, A4 => n10,
                           ZN => n44);
   U74 : INV_X1 port map( A => n34, ZN => n10);
   U75 : NOR2_X1 port map( A1 => tipo(0), A2 => n7, ZN => n45);
   U76 : XNOR2_X1 port map( A => n5, B => tipo(1), ZN => n49);
   U77 : INV_X1 port map( A => tipo(4), ZN => n9);
   U78 : INV_X1 port map( A => tipo(0), ZN => n5);
   U79 : INV_X1 port map( A => tipo(5), ZN => n11);

end SYN_Architectural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity logic_N32 is

   port( FUNC : in std_logic_vector (0 to 5);  DATA1, DATA2 : in 
         std_logic_vector (31 downto 0);  OUT_ALU : out std_logic_vector (31 
         downto 0));

end logic_N32;

architecture SYN_Architectural of logic_N32 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82,
      n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97
      , n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, 
      n110, n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, 
      n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, 
      n134, n135, n136, n137, n138, n139, n140, n1, n2, n3, n4, n5, n6, n7, n8,
      n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23,
      n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38
      , n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, 
      n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67
      , n68, n141, n142, n143, n144, n145, n146, n147, n148, n149, n150, n151, 
      n152, n153, n154, n155 : std_logic;

begin
   
   U173 : NAND3_X1 port map( A1 => n140, A2 => n154, A3 => FUNC(1), ZN => n136)
                           ;
   U2 : BUF_X1 port map( A => n71, Z => n12);
   U3 : BUF_X1 port map( A => n71, Z => n13);
   U4 : BUF_X1 port map( A => n71, Z => n14);
   U5 : BUF_X1 port map( A => n72, Z => n5);
   U6 : BUF_X1 port map( A => n72, Z => n4);
   U7 : BUF_X1 port map( A => n73, Z => n2);
   U8 : BUF_X1 port map( A => n73, Z => n1);
   U9 : BUF_X1 port map( A => n72, Z => n7);
   U10 : BUF_X1 port map( A => n72, Z => n8);
   U11 : OAI22_X1 port map( A1 => n86, A2 => n53, B1 => n87, B2 => n21, ZN => 
                           OUT_ALU(31));
   U12 : AOI21_X1 port map( B1 => n13, B2 => n53, A => n7, ZN => n87);
   U13 : AOI221_X1 port map( B1 => n12, B2 => n21, C1 => DATA1(31), C2 => n3, A
                           => n6, ZN => n86);
   U14 : INV_X1 port map( A => DATA2(31), ZN => n53);
   U15 : OAI22_X1 port map( A1 => n88, A2 => n54, B1 => n89, B2 => n22, ZN => 
                           OUT_ALU(30));
   U16 : AOI21_X1 port map( B1 => n13, B2 => n54, A => n7, ZN => n89);
   U17 : AOI221_X1 port map( B1 => n12, B2 => n22, C1 => DATA1(30), C2 => n2, A
                           => n6, ZN => n88);
   U18 : INV_X1 port map( A => DATA2(30), ZN => n54);
   U19 : OAI22_X1 port map( A1 => n92, A2 => n55, B1 => n93, B2 => n23, ZN => 
                           OUT_ALU(29));
   U20 : AOI21_X1 port map( B1 => n13, B2 => n55, A => n7, ZN => n93);
   U21 : AOI221_X1 port map( B1 => n12, B2 => n23, C1 => DATA1(29), C2 => n2, A
                           => n6, ZN => n92);
   U22 : INV_X1 port map( A => DATA2(29), ZN => n55);
   U23 : OAI22_X1 port map( A1 => n94, A2 => n56, B1 => n95, B2 => n24, ZN => 
                           OUT_ALU(28));
   U24 : AOI21_X1 port map( B1 => n13, B2 => n56, A => n7, ZN => n95);
   U25 : AOI221_X1 port map( B1 => n12, B2 => n24, C1 => DATA1(28), C2 => n2, A
                           => n6, ZN => n94);
   U26 : INV_X1 port map( A => DATA2(28), ZN => n56);
   U27 : OAI22_X1 port map( A1 => n96, A2 => n57, B1 => n97, B2 => n25, ZN => 
                           OUT_ALU(27));
   U28 : AOI21_X1 port map( B1 => n13, B2 => n57, A => n7, ZN => n97);
   U29 : AOI221_X1 port map( B1 => n12, B2 => n25, C1 => DATA1(27), C2 => n2, A
                           => n6, ZN => n96);
   U30 : INV_X1 port map( A => DATA2(27), ZN => n57);
   U31 : OAI22_X1 port map( A1 => n98, A2 => n58, B1 => n99, B2 => n26, ZN => 
                           OUT_ALU(26));
   U32 : AOI21_X1 port map( B1 => n13, B2 => n58, A => n7, ZN => n99);
   U33 : AOI221_X1 port map( B1 => n11, B2 => n26, C1 => DATA1(26), C2 => n2, A
                           => n5, ZN => n98);
   U34 : INV_X1 port map( A => DATA2(26), ZN => n58);
   U35 : OAI22_X1 port map( A1 => n100, A2 => n59, B1 => n101, B2 => n27, ZN =>
                           OUT_ALU(25));
   U36 : AOI21_X1 port map( B1 => n13, B2 => n59, A => n7, ZN => n101);
   U37 : AOI221_X1 port map( B1 => n12, B2 => n27, C1 => DATA1(25), C2 => n2, A
                           => n6, ZN => n100);
   U38 : INV_X1 port map( A => DATA2(25), ZN => n59);
   U39 : OAI22_X1 port map( A1 => n102, A2 => n60, B1 => n103, B2 => n28, ZN =>
                           OUT_ALU(24));
   U40 : AOI21_X1 port map( B1 => n14, B2 => n60, A => n7, ZN => n103);
   U41 : AOI221_X1 port map( B1 => n12, B2 => n28, C1 => DATA1(24), C2 => n2, A
                           => n6, ZN => n102);
   U42 : INV_X1 port map( A => DATA2(24), ZN => n60);
   U43 : OAI22_X1 port map( A1 => n104, A2 => n61, B1 => n105, B2 => n29, ZN =>
                           OUT_ALU(23));
   U44 : AOI21_X1 port map( B1 => n14, B2 => n61, A => n8, ZN => n105);
   U45 : AOI221_X1 port map( B1 => n11, B2 => n29, C1 => DATA1(23), C2 => n2, A
                           => n5, ZN => n104);
   U46 : INV_X1 port map( A => DATA2(23), ZN => n61);
   U47 : OAI22_X1 port map( A1 => n106, A2 => n62, B1 => n107, B2 => n30, ZN =>
                           OUT_ALU(22));
   U48 : AOI21_X1 port map( B1 => n14, B2 => n62, A => n8, ZN => n107);
   U49 : AOI221_X1 port map( B1 => n11, B2 => n30, C1 => DATA1(22), C2 => n2, A
                           => n5, ZN => n106);
   U50 : INV_X1 port map( A => DATA2(22), ZN => n62);
   U51 : OAI22_X1 port map( A1 => n108, A2 => n63, B1 => n109, B2 => n31, ZN =>
                           OUT_ALU(21));
   U52 : AOI21_X1 port map( B1 => n14, B2 => n63, A => n8, ZN => n109);
   U53 : AOI221_X1 port map( B1 => n11, B2 => n31, C1 => DATA1(21), C2 => n2, A
                           => n5, ZN => n108);
   U54 : INV_X1 port map( A => DATA2(21), ZN => n63);
   U55 : OAI22_X1 port map( A1 => n110, A2 => n64, B1 => n111, B2 => n32, ZN =>
                           OUT_ALU(20));
   U56 : AOI21_X1 port map( B1 => n14, B2 => n64, A => n8, ZN => n111);
   U57 : AOI221_X1 port map( B1 => n11, B2 => n32, C1 => DATA1(20), C2 => n2, A
                           => n5, ZN => n110);
   U58 : INV_X1 port map( A => DATA2(20), ZN => n64);
   U59 : OAI22_X1 port map( A1 => n114, A2 => n65, B1 => n115, B2 => n33, ZN =>
                           OUT_ALU(19));
   U60 : AOI21_X1 port map( B1 => n14, B2 => n65, A => n8, ZN => n115);
   U61 : AOI221_X1 port map( B1 => n11, B2 => n33, C1 => DATA1(19), C2 => n1, A
                           => n5, ZN => n114);
   U62 : INV_X1 port map( A => DATA2(19), ZN => n65);
   U63 : OAI22_X1 port map( A1 => n116, A2 => n66, B1 => n117, B2 => n34, ZN =>
                           OUT_ALU(18));
   U64 : AOI21_X1 port map( B1 => n14, B2 => n66, A => n8, ZN => n117);
   U65 : AOI221_X1 port map( B1 => n11, B2 => n34, C1 => DATA1(18), C2 => n1, A
                           => n5, ZN => n116);
   U66 : INV_X1 port map( A => DATA2(18), ZN => n66);
   U67 : OAI22_X1 port map( A1 => n118, A2 => n67, B1 => n119, B2 => n35, ZN =>
                           OUT_ALU(17));
   U68 : AOI21_X1 port map( B1 => n14, B2 => n67, A => n8, ZN => n119);
   U69 : AOI221_X1 port map( B1 => n11, B2 => n35, C1 => DATA1(17), C2 => n1, A
                           => n5, ZN => n118);
   U70 : INV_X1 port map( A => DATA2(17), ZN => n67);
   U71 : OAI22_X1 port map( A1 => n120, A2 => n68, B1 => n121, B2 => n36, ZN =>
                           OUT_ALU(16));
   U72 : AOI21_X1 port map( B1 => n14, B2 => n68, A => n8, ZN => n121);
   U73 : AOI221_X1 port map( B1 => n10, B2 => n36, C1 => DATA1(16), C2 => n1, A
                           => n4, ZN => n120);
   U74 : INV_X1 port map( A => DATA2(16), ZN => n68);
   U75 : OAI22_X1 port map( A1 => n122, A2 => n141, B1 => n123, B2 => n37, ZN 
                           => OUT_ALU(15));
   U76 : AOI21_X1 port map( B1 => n14, B2 => n141, A => n8, ZN => n123);
   U77 : AOI221_X1 port map( B1 => n10, B2 => n37, C1 => DATA1(15), C2 => n1, A
                           => n4, ZN => n122);
   U78 : INV_X1 port map( A => DATA2(15), ZN => n141);
   U79 : OAI22_X1 port map( A1 => n124, A2 => n142, B1 => n125, B2 => n38, ZN 
                           => OUT_ALU(14));
   U80 : AOI21_X1 port map( B1 => n14, B2 => n142, A => n8, ZN => n125);
   U81 : AOI221_X1 port map( B1 => n10, B2 => n38, C1 => DATA1(14), C2 => n1, A
                           => n4, ZN => n124);
   U82 : INV_X1 port map( A => DATA2(14), ZN => n142);
   U83 : OAI22_X1 port map( A1 => n126, A2 => n143, B1 => n127, B2 => n39, ZN 
                           => OUT_ALU(13));
   U84 : AOI21_X1 port map( B1 => n15, B2 => n143, A => n8, ZN => n127);
   U85 : AOI221_X1 port map( B1 => n10, B2 => n39, C1 => DATA1(13), C2 => n1, A
                           => n4, ZN => n126);
   U86 : INV_X1 port map( A => DATA2(13), ZN => n143);
   U87 : OAI22_X1 port map( A1 => n128, A2 => n144, B1 => n129, B2 => n40, ZN 
                           => OUT_ALU(12));
   U88 : AOI21_X1 port map( B1 => n15, B2 => n144, A => n8, ZN => n129);
   U89 : AOI221_X1 port map( B1 => n10, B2 => n40, C1 => DATA1(12), C2 => n1, A
                           => n4, ZN => n128);
   U90 : INV_X1 port map( A => DATA2(12), ZN => n144);
   U91 : OAI22_X1 port map( A1 => n130, A2 => n145, B1 => n131, B2 => n41, ZN 
                           => OUT_ALU(11));
   U92 : AOI21_X1 port map( B1 => n15, B2 => n145, A => n9, ZN => n131);
   U93 : AOI221_X1 port map( B1 => n10, B2 => n41, C1 => DATA1(11), C2 => n1, A
                           => n4, ZN => n130);
   U94 : INV_X1 port map( A => DATA2(11), ZN => n145);
   U95 : OAI22_X1 port map( A1 => n132, A2 => n146, B1 => n133, B2 => n42, ZN 
                           => OUT_ALU(10));
   U96 : AOI21_X1 port map( B1 => n15, B2 => n146, A => n9, ZN => n133);
   U97 : AOI221_X1 port map( B1 => n10, B2 => n42, C1 => DATA1(10), C2 => n1, A
                           => n4, ZN => n132);
   U98 : INV_X1 port map( A => DATA2(10), ZN => n146);
   U99 : OAI22_X1 port map( A1 => n69, A2 => n147, B1 => n70, B2 => n43, ZN => 
                           OUT_ALU(9));
   U100 : AOI21_X1 port map( B1 => n13, B2 => n147, A => n7, ZN => n70);
   U101 : AOI221_X1 port map( B1 => n10, B2 => n43, C1 => n3, C2 => DATA1(9), A
                           => n4, ZN => n69);
   U102 : INV_X1 port map( A => DATA2(9), ZN => n147);
   U103 : OAI22_X1 port map( A1 => n74, A2 => n148, B1 => n75, B2 => n44, ZN =>
                           OUT_ALU(8));
   U104 : AOI21_X1 port map( B1 => n12, B2 => n148, A => n6, ZN => n75);
   U105 : AOI221_X1 port map( B1 => n10, B2 => n44, C1 => DATA1(8), C2 => n3, A
                           => n4, ZN => n74);
   U106 : INV_X1 port map( A => DATA2(8), ZN => n148);
   U107 : OAI22_X1 port map( A1 => n76, A2 => n149, B1 => n77, B2 => n45, ZN =>
                           OUT_ALU(7));
   U108 : AOI21_X1 port map( B1 => n13, B2 => n149, A => n7, ZN => n77);
   U109 : AOI221_X1 port map( B1 => n10, B2 => n45, C1 => DATA1(7), C2 => n3, A
                           => n4, ZN => n76);
   U110 : INV_X1 port map( A => DATA2(7), ZN => n149);
   U111 : OAI22_X1 port map( A1 => n78, A2 => n150, B1 => n79, B2 => n46, ZN =>
                           OUT_ALU(6));
   U112 : AOI21_X1 port map( B1 => n12, B2 => n150, A => n6, ZN => n79);
   U113 : AOI221_X1 port map( B1 => n10, B2 => n46, C1 => DATA1(6), C2 => n3, A
                           => n4, ZN => n78);
   U114 : INV_X1 port map( A => DATA2(6), ZN => n150);
   U115 : OAI22_X1 port map( A1 => n80, A2 => n151, B1 => n81, B2 => n47, ZN =>
                           OUT_ALU(5));
   U116 : AOI21_X1 port map( B1 => n12, B2 => n151, A => n6, ZN => n81);
   U117 : AOI221_X1 port map( B1 => n11, B2 => n47, C1 => DATA1(5), C2 => n3, A
                           => n5, ZN => n80);
   U118 : INV_X1 port map( A => DATA2(5), ZN => n151);
   U119 : OAI22_X1 port map( A1 => n82, A2 => n20, B1 => n83, B2 => n48, ZN => 
                           OUT_ALU(4));
   U120 : AOI21_X1 port map( B1 => n13, B2 => n20, A => n7, ZN => n83);
   U121 : AOI221_X1 port map( B1 => n11, B2 => n48, C1 => DATA1(4), C2 => n3, A
                           => n5, ZN => n82);
   U122 : OAI22_X1 port map( A1 => n84, A2 => n19, B1 => n85, B2 => n49, ZN => 
                           OUT_ALU(3));
   U123 : AOI21_X1 port map( B1 => n13, B2 => n19, A => n7, ZN => n85);
   U124 : AOI221_X1 port map( B1 => n11, B2 => n49, C1 => DATA1(3), C2 => n3, A
                           => n5, ZN => n84);
   U125 : OAI22_X1 port map( A1 => n90, A2 => n18, B1 => n91, B2 => n50, ZN => 
                           OUT_ALU(2));
   U126 : AOI21_X1 port map( B1 => n13, B2 => n18, A => n7, ZN => n91);
   U127 : AOI221_X1 port map( B1 => n12, B2 => n50, C1 => DATA1(2), C2 => n2, A
                           => n6, ZN => n90);
   U128 : OAI22_X1 port map( A1 => n112, A2 => n17, B1 => n113, B2 => n51, ZN 
                           => OUT_ALU(1));
   U129 : AOI21_X1 port map( B1 => n14, B2 => n17, A => n8, ZN => n113);
   U130 : AOI221_X1 port map( B1 => n11, B2 => n51, C1 => DATA1(1), C2 => n1, A
                           => n5, ZN => n112);
   U131 : OAI22_X1 port map( A1 => n134, A2 => n16, B1 => n135, B2 => n52, ZN 
                           => OUT_ALU(0));
   U132 : AOI21_X1 port map( B1 => n12, B2 => n16, A => n6, ZN => n135);
   U133 : AOI221_X1 port map( B1 => n10, B2 => n52, C1 => DATA1(0), C2 => n1, A
                           => n4, ZN => n134);
   U134 : BUF_X1 port map( A => n72, Z => n6);
   U135 : BUF_X1 port map( A => n71, Z => n11);
   U136 : BUF_X1 port map( A => n71, Z => n10);
   U137 : BUF_X1 port map( A => n73, Z => n3);
   U138 : INV_X1 port map( A => DATA1(12), ZN => n40);
   U139 : INV_X1 port map( A => DATA1(23), ZN => n29);
   U140 : INV_X1 port map( A => DATA1(14), ZN => n38);
   U141 : INV_X1 port map( A => DATA1(17), ZN => n35);
   U142 : INV_X1 port map( A => DATA1(21), ZN => n31);
   U143 : INV_X1 port map( A => DATA1(13), ZN => n39);
   U144 : INV_X1 port map( A => DATA1(22), ZN => n30);
   U145 : INV_X1 port map( A => DATA1(16), ZN => n36);
   U146 : INV_X1 port map( A => DATA1(15), ZN => n37);
   U147 : INV_X1 port map( A => DATA1(9), ZN => n43);
   U148 : INV_X1 port map( A => DATA1(11), ZN => n41);
   U149 : INV_X1 port map( A => DATA1(10), ZN => n42);
   U150 : INV_X1 port map( A => DATA1(8), ZN => n44);
   U151 : INV_X1 port map( A => DATA1(7), ZN => n45);
   U152 : INV_X1 port map( A => DATA1(2), ZN => n50);
   U153 : INV_X1 port map( A => DATA1(3), ZN => n49);
   U154 : INV_X1 port map( A => DATA1(28), ZN => n24);
   U155 : INV_X1 port map( A => DATA1(27), ZN => n25);
   U156 : INV_X1 port map( A => DATA1(26), ZN => n26);
   U157 : INV_X1 port map( A => DATA1(25), ZN => n27);
   U158 : INV_X1 port map( A => DATA1(24), ZN => n28);
   U159 : INV_X1 port map( A => DATA1(18), ZN => n34);
   U160 : INV_X1 port map( A => DATA1(0), ZN => n52);
   U161 : INV_X1 port map( A => DATA1(29), ZN => n23);
   U162 : INV_X1 port map( A => DATA1(4), ZN => n48);
   U163 : INV_X1 port map( A => DATA1(6), ZN => n46);
   U164 : INV_X1 port map( A => DATA1(31), ZN => n21);
   U165 : INV_X1 port map( A => DATA1(19), ZN => n33);
   U166 : INV_X1 port map( A => DATA1(20), ZN => n32);
   U167 : INV_X1 port map( A => DATA1(1), ZN => n51);
   U168 : INV_X1 port map( A => DATA1(5), ZN => n47);
   U169 : INV_X1 port map( A => DATA1(30), ZN => n22);
   U170 : OAI21_X1 port map( B1 => FUNC(5), B2 => n136, A => n137, ZN => n72);
   U171 : OR3_X1 port map( A1 => n138, A2 => FUNC(2), A3 => n155, ZN => n137);
   U172 : NAND4_X1 port map( A1 => FUNC(3), A2 => FUNC(4), A3 => n153, A4 => 
                           n152, ZN => n138);
   U174 : INV_X1 port map( A => FUNC(0), ZN => n152);
   U175 : NOR3_X1 port map( A1 => FUNC(3), A2 => FUNC(0), A3 => FUNC(4), ZN => 
                           n140);
   U176 : AOI21_X1 port map( B1 => n155, B2 => FUNC(2), A => n138, ZN => n73);
   U177 : INV_X1 port map( A => FUNC(2), ZN => n154);
   U178 : NAND2_X1 port map( A1 => n136, A2 => n139, ZN => n71);
   U179 : NAND4_X1 port map( A1 => FUNC(2), A2 => n140, A3 => n155, A4 => n153,
                           ZN => n139);
   U180 : INV_X1 port map( A => FUNC(5), ZN => n155);
   U181 : INV_X1 port map( A => FUNC(1), ZN => n153);
   U182 : CLKBUF_X1 port map( A => n72, Z => n9);
   U183 : CLKBUF_X1 port map( A => n71, Z => n15);
   U184 : INV_X1 port map( A => DATA2(0), ZN => n16);
   U185 : INV_X1 port map( A => DATA2(1), ZN => n17);
   U186 : INV_X1 port map( A => DATA2(2), ZN => n18);
   U187 : INV_X1 port map( A => DATA2(3), ZN => n19);
   U188 : INV_X1 port map( A => DATA2(4), ZN => n20);

end SYN_Architectural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity sign_eval_N_in26_N_out32 is

   port( IR_out : in std_logic_vector (25 downto 0);  signed_val : in std_logic
         ;  Immediate : out std_logic_vector (31 downto 0));

end sign_eval_N_in26_N_out32;

architecture SYN_BHV of sign_eval_N_in26_N_out32 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal N0, n1 : std_logic;

begin
   Immediate <= ( N0, N0, N0, N0, N0, N0, IR_out(25), IR_out(24), IR_out(23), 
      IR_out(22), IR_out(21), IR_out(20), IR_out(19), IR_out(18), IR_out(17), 
      IR_out(16), IR_out(15), IR_out(14), IR_out(13), IR_out(12), IR_out(11), 
      IR_out(10), IR_out(9), IR_out(8), IR_out(7), IR_out(6), IR_out(5), 
      IR_out(4), IR_out(3), IR_out(2), IR_out(1), IR_out(0) );
   
   U1 : NOR2_X1 port map( A1 => signed_val, A2 => n1, ZN => N0);
   U2 : INV_X1 port map( A => IR_out(25), ZN => n1);

end SYN_BHV;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity sign_eval_N_in16_N_out32 is

   port( IR_out : in std_logic_vector (15 downto 0);  signed_val : in std_logic
         ;  Immediate : out std_logic_vector (31 downto 0));

end sign_eval_N_in16_N_out32;

architecture SYN_BHV of sign_eval_N_in16_N_out32 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal N0, n1 : std_logic;

begin
   Immediate <= ( N0, N0, N0, N0, N0, N0, N0, N0, N0, N0, N0, N0, N0, N0, N0, 
      N0, IR_out(15), IR_out(14), IR_out(13), IR_out(12), IR_out(11), 
      IR_out(10), IR_out(9), IR_out(8), IR_out(7), IR_out(6), IR_out(5), 
      IR_out(4), IR_out(3), IR_out(2), IR_out(1), IR_out(0) );
   
   U1 : NOR2_X1 port map( A1 => signed_val, A2 => n1, ZN => N0);
   U2 : INV_X1 port map( A => IR_out(15), ZN => n1);

end SYN_BHV;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity sign_eval_N_in5_N_out32 is

   port( IR_out : in std_logic_vector (4 downto 0);  signed_val : in std_logic;
         Immediate : out std_logic_vector (31 downto 0));

end sign_eval_N_in5_N_out32;

architecture SYN_BHV of sign_eval_N_in5_N_out32 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal N0, n1 : std_logic;

begin
   Immediate <= ( N0, N0, N0, N0, N0, N0, N0, N0, N0, N0, N0, N0, N0, N0, N0, 
      N0, N0, N0, N0, N0, N0, N0, N0, N0, N0, N0, N0, IR_out(4), IR_out(3), 
      IR_out(2), IR_out(1), IR_out(0) );
   
   U1 : NOR2_X1 port map( A1 => signed_val, A2 => n1, ZN => N0);
   U2 : INV_X1 port map( A => IR_out(4), ZN => n1);

end SYN_BHV;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_0 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_0;

architecture SYN_STRUCTURAL of MUX21_0 is

   component ND2_766
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_767
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component ND2_0
      port( A, B : in std_logic;  Y : out std_logic);
   end component;
   
   component IV_0
      port( A : in std_logic;  Y : out std_logic);
   end component;
   
   signal SB, Y1, Y2 : std_logic;

begin
   
   UIV : IV_0 port map( A => S, Y => SB);
   UND1 : ND2_0 port map( A => A, B => S, Y => Y1);
   UND2 : ND2_767 port map( A => B, B => SB, Y => Y2);
   UND3 : ND2_766 port map( A => Y1, B => Y2, Y => Y);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity load_data is

   port( data_in : in std_logic_vector (31 downto 0);  signed_val, load_op : in
         std_logic;  load_type : in std_logic_vector (1 downto 0);  data_out : 
         out std_logic_vector (31 downto 0));

end load_data;

architecture SYN_bhv_load of load_data is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N36, N37, N38, N39, N40, N41, N42, N43, N44, N45, N46, N47, N48, N49,
      N50, N51, N52, N53, N54, N55, N56, N57, N58, N59, N60, N61, N62, N63, N64
      , N65, N66, N67, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, 
      n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30
      , n1, n2, n3, n31, n32 : std_logic;

begin
   
   data_out_reg_31_inst : DLH_X1 port map( G => load_op, D => N67, Q => 
                           data_out(31));
   data_out_reg_30_inst : DLH_X1 port map( G => load_op, D => N66, Q => 
                           data_out(30));
   data_out_reg_29_inst : DLH_X1 port map( G => load_op, D => N65, Q => 
                           data_out(29));
   data_out_reg_28_inst : DLH_X1 port map( G => load_op, D => N64, Q => 
                           data_out(28));
   data_out_reg_27_inst : DLH_X1 port map( G => load_op, D => N63, Q => 
                           data_out(27));
   data_out_reg_26_inst : DLH_X1 port map( G => load_op, D => N62, Q => 
                           data_out(26));
   data_out_reg_25_inst : DLH_X1 port map( G => load_op, D => N61, Q => 
                           data_out(25));
   data_out_reg_24_inst : DLH_X1 port map( G => load_op, D => N60, Q => 
                           data_out(24));
   data_out_reg_23_inst : DLH_X1 port map( G => load_op, D => N59, Q => 
                           data_out(23));
   data_out_reg_22_inst : DLH_X1 port map( G => load_op, D => N58, Q => 
                           data_out(22));
   data_out_reg_21_inst : DLH_X1 port map( G => load_op, D => N57, Q => 
                           data_out(21));
   data_out_reg_20_inst : DLH_X1 port map( G => load_op, D => N56, Q => 
                           data_out(20));
   data_out_reg_19_inst : DLH_X1 port map( G => load_op, D => N55, Q => 
                           data_out(19));
   data_out_reg_18_inst : DLH_X1 port map( G => load_op, D => N54, Q => 
                           data_out(18));
   data_out_reg_17_inst : DLH_X1 port map( G => load_op, D => N53, Q => 
                           data_out(17));
   data_out_reg_16_inst : DLH_X1 port map( G => load_op, D => N52, Q => 
                           data_out(16));
   data_out_reg_15_inst : DLH_X1 port map( G => load_op, D => N51, Q => 
                           data_out(15));
   data_out_reg_14_inst : DLH_X1 port map( G => load_op, D => N50, Q => 
                           data_out(14));
   data_out_reg_13_inst : DLH_X1 port map( G => load_op, D => N49, Q => 
                           data_out(13));
   data_out_reg_12_inst : DLH_X1 port map( G => load_op, D => N48, Q => 
                           data_out(12));
   data_out_reg_11_inst : DLH_X1 port map( G => load_op, D => N47, Q => 
                           data_out(11));
   data_out_reg_10_inst : DLH_X1 port map( G => load_op, D => N46, Q => 
                           data_out(10));
   data_out_reg_9_inst : DLH_X1 port map( G => load_op, D => N45, Q => 
                           data_out(9));
   data_out_reg_8_inst : DLH_X1 port map( G => load_op, D => N44, Q => 
                           data_out(8));
   data_out_reg_7_inst : DLH_X1 port map( G => load_op, D => N43, Q => 
                           data_out(7));
   data_out_reg_6_inst : DLH_X1 port map( G => load_op, D => N42, Q => 
                           data_out(6));
   data_out_reg_5_inst : DLH_X1 port map( G => load_op, D => N41, Q => 
                           data_out(5));
   data_out_reg_4_inst : DLH_X1 port map( G => load_op, D => N40, Q => 
                           data_out(4));
   data_out_reg_3_inst : DLH_X1 port map( G => load_op, D => N39, Q => 
                           data_out(3));
   data_out_reg_2_inst : DLH_X1 port map( G => load_op, D => N38, Q => 
                           data_out(2));
   data_out_reg_1_inst : DLH_X1 port map( G => load_op, D => N37, Q => 
                           data_out(1));
   data_out_reg_0_inst : DLH_X1 port map( G => load_op, D => N36, Q => 
                           data_out(0));
   U2 : INV_X1 port map( A => n4, ZN => n3);
   U3 : BUF_X1 port map( A => n5, Z => n1);
   U4 : BUF_X1 port map( A => n5, Z => n2);
   U5 : OAI21_X1 port map( B1 => n4, B2 => n32, A => n1, ZN => N67);
   U6 : NAND2_X1 port map( A1 => load_type(1), A2 => load_type(0), ZN => n4);
   U7 : NAND2_X1 port map( A1 => n31, A2 => n29, ZN => n30);
   U8 : INV_X1 port map( A => load_type(0), ZN => n31);
   U9 : OR2_X1 port map( A1 => load_type(1), A2 => load_type(0), ZN => n29);
   U10 : OR3_X1 port map( A1 => signed_val, A2 => n32, A3 => n29, ZN => n5);
   U11 : INV_X1 port map( A => data_in(31), ZN => n32);
   U12 : NAND2_X1 port map( A1 => n2, A2 => n28, ZN => N44);
   U13 : NAND2_X1 port map( A1 => data_in(8), A2 => load_type(0), ZN => n28);
   U14 : NAND2_X1 port map( A1 => n2, A2 => n27, ZN => N45);
   U15 : NAND2_X1 port map( A1 => data_in(9), A2 => load_type(0), ZN => n27);
   U16 : NAND2_X1 port map( A1 => n2, A2 => n26, ZN => N46);
   U17 : NAND2_X1 port map( A1 => data_in(10), A2 => load_type(0), ZN => n26);
   U18 : NAND2_X1 port map( A1 => n2, A2 => n25, ZN => N47);
   U19 : NAND2_X1 port map( A1 => data_in(11), A2 => load_type(0), ZN => n25);
   U20 : NAND2_X1 port map( A1 => n2, A2 => n24, ZN => N48);
   U21 : NAND2_X1 port map( A1 => data_in(12), A2 => load_type(0), ZN => n24);
   U22 : NAND2_X1 port map( A1 => n2, A2 => n23, ZN => N49);
   U23 : NAND2_X1 port map( A1 => data_in(13), A2 => load_type(0), ZN => n23);
   U24 : NAND2_X1 port map( A1 => n2, A2 => n22, ZN => N50);
   U25 : NAND2_X1 port map( A1 => data_in(14), A2 => load_type(0), ZN => n22);
   U26 : NAND2_X1 port map( A1 => n2, A2 => n21, ZN => N51);
   U27 : NAND2_X1 port map( A1 => data_in(15), A2 => load_type(0), ZN => n21);
   U28 : NAND2_X1 port map( A1 => n1, A2 => n16, ZN => N56);
   U29 : NAND2_X1 port map( A1 => data_in(20), A2 => n3, ZN => n16);
   U30 : NAND2_X1 port map( A1 => n1, A2 => n15, ZN => N57);
   U31 : NAND2_X1 port map( A1 => data_in(21), A2 => n3, ZN => n15);
   U32 : NAND2_X1 port map( A1 => n1, A2 => n14, ZN => N58);
   U33 : NAND2_X1 port map( A1 => data_in(22), A2 => n3, ZN => n14);
   U34 : NAND2_X1 port map( A1 => n1, A2 => n13, ZN => N59);
   U35 : NAND2_X1 port map( A1 => data_in(23), A2 => n3, ZN => n13);
   U36 : NAND2_X1 port map( A1 => n1, A2 => n12, ZN => N60);
   U37 : NAND2_X1 port map( A1 => data_in(24), A2 => n3, ZN => n12);
   U38 : NAND2_X1 port map( A1 => n1, A2 => n11, ZN => N61);
   U39 : NAND2_X1 port map( A1 => data_in(25), A2 => n3, ZN => n11);
   U40 : NAND2_X1 port map( A1 => n1, A2 => n10, ZN => N62);
   U41 : NAND2_X1 port map( A1 => data_in(26), A2 => n3, ZN => n10);
   U42 : NAND2_X1 port map( A1 => n1, A2 => n9, ZN => N63);
   U43 : NAND2_X1 port map( A1 => data_in(27), A2 => n3, ZN => n9);
   U44 : NAND2_X1 port map( A1 => n1, A2 => n8, ZN => N64);
   U45 : NAND2_X1 port map( A1 => data_in(28), A2 => n3, ZN => n8);
   U46 : NAND2_X1 port map( A1 => n1, A2 => n7, ZN => N65);
   U47 : NAND2_X1 port map( A1 => data_in(29), A2 => n3, ZN => n7);
   U48 : NAND2_X1 port map( A1 => n1, A2 => n6, ZN => N66);
   U49 : NAND2_X1 port map( A1 => data_in(30), A2 => n3, ZN => n6);
   U50 : NAND2_X1 port map( A1 => n2, A2 => n20, ZN => N52);
   U51 : NAND2_X1 port map( A1 => data_in(16), A2 => n3, ZN => n20);
   U52 : NAND2_X1 port map( A1 => n2, A2 => n19, ZN => N53);
   U53 : NAND2_X1 port map( A1 => data_in(17), A2 => n3, ZN => n19);
   U54 : NAND2_X1 port map( A1 => n2, A2 => n18, ZN => N54);
   U55 : NAND2_X1 port map( A1 => data_in(18), A2 => n3, ZN => n18);
   U56 : NAND2_X1 port map( A1 => n2, A2 => n17, ZN => N55);
   U57 : NAND2_X1 port map( A1 => data_in(19), A2 => n3, ZN => n17);
   U58 : AND2_X1 port map( A1 => data_in(0), A2 => n30, ZN => N36);
   U59 : AND2_X1 port map( A1 => data_in(1), A2 => n30, ZN => N37);
   U60 : AND2_X1 port map( A1 => data_in(2), A2 => n30, ZN => N38);
   U61 : AND2_X1 port map( A1 => data_in(3), A2 => n30, ZN => N39);
   U62 : AND2_X1 port map( A1 => data_in(4), A2 => n30, ZN => N40);
   U63 : AND2_X1 port map( A1 => data_in(5), A2 => n30, ZN => N41);
   U64 : AND2_X1 port map( A1 => data_in(6), A2 => n30, ZN => N42);
   U65 : AND2_X1 port map( A1 => data_in(7), A2 => n30, ZN => N43);

end SYN_bhv_load;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity COND_BT_NBIT32 is

   port( ZERO_BIT, OPCODE_0, branch_op : in std_logic;  con_sign : out 
         std_logic);

end COND_BT_NBIT32;

architecture SYN_BHV of COND_BT_NBIT32 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ZERO_BIT, B => OPCODE_0, Z => n1);
   U2 : AND2_X1 port map( A1 => branch_op, A2 => n1, ZN => con_sign);

end SYN_BHV;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity zero_eval_NBIT32 is

   port( input : in std_logic_vector (31 downto 0);  res : out std_logic);

end zero_eval_NBIT32;

architecture SYN_bhv of zero_eval_NBIT32 is

   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10 : std_logic;

begin
   
   U1 : NOR4_X1 port map( A1 => input(23), A2 => input(22), A3 => input(21), A4
                           => input(20), ZN => n6);
   U2 : NOR4_X1 port map( A1 => input(9), A2 => input(8), A3 => input(7), A4 =>
                           input(6), ZN => n10);
   U3 : NOR4_X1 port map( A1 => input(5), A2 => input(4), A3 => input(3), A4 =>
                           input(31), ZN => n9);
   U4 : NOR4_X1 port map( A1 => input(30), A2 => input(2), A3 => input(29), A4 
                           => input(28), ZN => n8);
   U5 : NOR4_X1 port map( A1 => input(27), A2 => input(26), A3 => input(25), A4
                           => input(24), ZN => n7);
   U6 : NAND4_X1 port map( A1 => n3, A2 => n4, A3 => n5, A4 => n6, ZN => n2);
   U7 : NOR4_X1 port map( A1 => input(12), A2 => input(11), A3 => input(10), A4
                           => input(0), ZN => n3);
   U8 : NOR4_X1 port map( A1 => input(16), A2 => input(15), A3 => input(14), A4
                           => input(13), ZN => n4);
   U9 : NOR4_X1 port map( A1 => input(1), A2 => input(19), A3 => input(18), A4 
                           => input(17), ZN => n5);
   U10 : NOR2_X1 port map( A1 => n1, A2 => n2, ZN => res);
   U11 : NAND4_X1 port map( A1 => n7, A2 => n8, A3 => n9, A4 => n10, ZN => n1);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ALU_N32 is

   port( CLK : in std_logic;  FUNC : in std_logic_vector (0 to 5);  DATA1, 
         DATA2 : in std_logic_vector (31 downto 0);  OUT_ALU : out 
         std_logic_vector (31 downto 0));

end ALU_N32;

architecture SYN_Architectural of ALU_N32 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component P4_ADDER_NBIT32
      port( A, B : in std_logic_vector (31 downto 0);  Cin : in std_logic;  S :
            out std_logic_vector (31 downto 0);  Cout : out std_logic);
   end component;
   
   component SHIFTER_GENERIC_N32
      port( A : in std_logic_vector (31 downto 0);  B : in std_logic_vector (4 
            downto 0);  LOGIC_ARITH, LEFT_RIGHT, SHIFT_ROTATE : in std_logic;  
            OUTPUT : out std_logic_vector (31 downto 0));
   end component;
   
   component comparator
      port( DATA1 : in std_logic_vector (31 downto 0);  DATA2i : in std_logic; 
            tipo : in std_logic_vector (0 to 5);  OUTALU : out std_logic_vector
            (31 downto 0));
   end component;
   
   component logic_N32
      port( FUNC : in std_logic_vector (0 to 5);  DATA1, DATA2 : in 
            std_logic_vector (31 downto 0);  OUT_ALU : out std_logic_vector (31
            downto 0));
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal OUTPUT_alu_i_31_port, OUTPUT_alu_i_30_port, OUTPUT_alu_i_29_port, 
      OUTPUT_alu_i_28_port, OUTPUT_alu_i_27_port, OUTPUT_alu_i_26_port, 
      OUTPUT_alu_i_25_port, OUTPUT_alu_i_24_port, OUTPUT_alu_i_23_port, 
      OUTPUT_alu_i_22_port, OUTPUT_alu_i_21_port, OUTPUT_alu_i_20_port, 
      OUTPUT_alu_i_19_port, OUTPUT_alu_i_18_port, OUTPUT_alu_i_17_port, 
      OUTPUT_alu_i_16_port, OUTPUT_alu_i_15_port, OUTPUT_alu_i_14_port, 
      OUTPUT_alu_i_13_port, OUTPUT_alu_i_12_port, OUTPUT_alu_i_11_port, 
      OUTPUT_alu_i_10_port, OUTPUT_alu_i_9_port, OUTPUT_alu_i_8_port, 
      OUTPUT_alu_i_7_port, OUTPUT_alu_i_6_port, OUTPUT_alu_i_5_port, 
      OUTPUT_alu_i_4_port, OUTPUT_alu_i_3_port, OUTPUT_alu_i_2_port, 
      OUTPUT_alu_i_1_port, OUTPUT_alu_i_0_port, OUTPUT4_31_port, 
      OUTPUT4_30_port, OUTPUT4_29_port, OUTPUT4_28_port, OUTPUT4_27_port, 
      OUTPUT4_26_port, OUTPUT4_25_port, OUTPUT4_24_port, OUTPUT4_23_port, 
      OUTPUT4_22_port, OUTPUT4_21_port, OUTPUT4_20_port, OUTPUT4_19_port, 
      OUTPUT4_18_port, OUTPUT4_17_port, OUTPUT4_16_port, OUTPUT4_15_port, 
      OUTPUT4_14_port, OUTPUT4_13_port, OUTPUT4_12_port, OUTPUT4_11_port, 
      OUTPUT4_10_port, OUTPUT4_9_port, OUTPUT4_8_port, OUTPUT4_7_port, 
      OUTPUT4_6_port, OUTPUT4_5_port, OUTPUT4_4_port, OUTPUT4_3_port, 
      OUTPUT4_2_port, OUTPUT4_1_port, OUTPUT4_0_port, OUTPUT2_31_port, 
      OUTPUT2_30_port, OUTPUT2_29_port, OUTPUT2_28_port, OUTPUT2_27_port, 
      OUTPUT2_26_port, OUTPUT2_25_port, OUTPUT2_24_port, OUTPUT2_23_port, 
      OUTPUT2_22_port, OUTPUT2_21_port, OUTPUT2_20_port, OUTPUT2_19_port, 
      OUTPUT2_18_port, OUTPUT2_17_port, OUTPUT2_16_port, OUTPUT2_15_port, 
      OUTPUT2_14_port, OUTPUT2_13_port, OUTPUT2_12_port, OUTPUT2_11_port, 
      OUTPUT2_10_port, OUTPUT2_9_port, OUTPUT2_8_port, OUTPUT2_7_port, 
      OUTPUT2_6_port, OUTPUT2_5_port, OUTPUT2_4_port, OUTPUT2_3_port, 
      OUTPUT2_2_port, OUTPUT2_1_port, OUTPUT2_0_port, Cout_i, OUTPUT3_0_port, 
      LOGIC_ARITH_i, LEFT_RIGHT_i, SHIFT_ROTATE_i, OUTPUT1_31_port, 
      OUTPUT1_30_port, OUTPUT1_29_port, OUTPUT1_28_port, OUTPUT1_27_port, 
      OUTPUT1_26_port, OUTPUT1_25_port, OUTPUT1_24_port, OUTPUT1_23_port, 
      OUTPUT1_22_port, OUTPUT1_21_port, OUTPUT1_20_port, OUTPUT1_19_port, 
      OUTPUT1_18_port, OUTPUT1_17_port, OUTPUT1_16_port, OUTPUT1_15_port, 
      OUTPUT1_14_port, OUTPUT1_13_port, OUTPUT1_12_port, OUTPUT1_11_port, 
      OUTPUT1_10_port, OUTPUT1_9_port, OUTPUT1_8_port, OUTPUT1_7_port, 
      OUTPUT1_6_port, OUTPUT1_5_port, OUTPUT1_4_port, OUTPUT1_3_port, 
      OUTPUT1_2_port, OUTPUT1_1_port, OUTPUT1_0_port, data1i_31_port, 
      data1i_30_port, data1i_29_port, data1i_28_port, data1i_27_port, 
      data1i_26_port, data1i_25_port, data1i_24_port, data1i_23_port, 
      data1i_22_port, data1i_21_port, data1i_20_port, data1i_19_port, 
      data1i_18_port, data1i_17_port, data1i_16_port, data1i_15_port, 
      data1i_14_port, data1i_13_port, data1i_12_port, data1i_11_port, 
      data1i_10_port, data1i_9_port, data1i_8_port, data1i_7_port, 
      data1i_6_port, data1i_5_port, data1i_4_port, data1i_3_port, data1i_2_port
      , data1i_1_port, data1i_0_port, data2i_31_port, data2i_30_port, 
      data2i_29_port, data2i_28_port, data2i_27_port, data2i_26_port, 
      data2i_25_port, data2i_24_port, data2i_23_port, data2i_22_port, 
      data2i_21_port, data2i_20_port, data2i_19_port, data2i_18_port, 
      data2i_17_port, data2i_16_port, data2i_15_port, data2i_14_port, 
      data2i_13_port, data2i_12_port, data2i_11_port, data2i_10_port, 
      data2i_9_port, data2i_8_port, data2i_7_port, data2i_6_port, data2i_5_port
      , data2i_4_port, data2i_3_port, data2i_2_port, data2i_1_port, 
      data2i_0_port, Cin_i, N139, N141, N142, N143, N144, N145, N146, N147, 
      N148, N149, N150, N151, N152, N153, N154, N155, N156, N157, N158, N159, 
      N160, N161, N162, N163, N164, N165, N166, N167, N168, N169, N170, N171, 
      N172, N173, N174, N175, N176, N177, N178, N179, N180, N181, N182, N183, 
      N184, N185, N186, N187, N188, N189, N190, N191, N192, N193, N194, N195, 
      N196, N197, N198, N199, N200, N201, N202, N203, N204, N205, N206, n48, 
      n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64
      , n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, 
      n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93
      , n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106,
      n107, n108, n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, 
      n119, n120, n121, n122, n123, n124, n125, n126, n127, n128, n129, n130, 
      n131, n132, n133, n134, n135, n136, n137, n138, n139_port, n140, 
      n141_port, n142_port, n143_port, n144_port, n145_port, n146_port, 
      n147_port, n148_port, n149_port, n150_port, n151_port, n152_port, 
      n153_port, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, 
      n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29
      , n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, 
      n44, n45, n46, n47, n49, n154_port, n155_port, n156_port, n157_port, 
      n158_port, n159_port, n160_port, n161_port, n162_port, n163_port, 
      n164_port, n165_port, n166_port, n167_port, n168_port, n169_port, 
      n170_port, n171_port, n172_port, n173_port, n174_port, n_1089, n_1090, 
      n_1091, n_1092, n_1093, n_1094, n_1095, n_1096, n_1097, n_1098, n_1099, 
      n_1100, n_1101, n_1102, n_1103, n_1104, n_1105, n_1106, n_1107, n_1108, 
      n_1109, n_1110, n_1111, n_1112, n_1113, n_1114, n_1115, n_1116, n_1117, 
      n_1118, n_1119, n_1120, n_1121, n_1122, n_1123, n_1124, n_1125, n_1126, 
      n_1127, n_1128, n_1129, n_1130, n_1131, n_1132, n_1133, n_1134, n_1135, 
      n_1136, n_1137, n_1138, n_1139, n_1140, n_1141, n_1142, n_1143, n_1144, 
      n_1145, n_1146, n_1147, n_1148, n_1149, n_1150, n_1151 : std_logic;

begin
   
   Cin_i_reg : DLH_X1 port map( G => n19, D => n1, Q => Cin_i);
   data2i_reg_31_inst : DLH_X1 port map( G => n19, D => N205, Q => 
                           data2i_31_port);
   data2i_reg_30_inst : DLH_X1 port map( G => n19, D => N204, Q => 
                           data2i_30_port);
   data2i_reg_29_inst : DLH_X1 port map( G => n19, D => N203, Q => 
                           data2i_29_port);
   data2i_reg_28_inst : DLH_X1 port map( G => n19, D => N202, Q => 
                           data2i_28_port);
   data2i_reg_27_inst : DLH_X1 port map( G => n19, D => N201, Q => 
                           data2i_27_port);
   data2i_reg_26_inst : DLH_X1 port map( G => n19, D => N200, Q => 
                           data2i_26_port);
   data2i_reg_25_inst : DLH_X1 port map( G => n19, D => N199, Q => 
                           data2i_25_port);
   data2i_reg_24_inst : DLH_X1 port map( G => n19, D => N198, Q => 
                           data2i_24_port);
   data2i_reg_23_inst : DLH_X1 port map( G => n19, D => N197, Q => 
                           data2i_23_port);
   data2i_reg_22_inst : DLH_X1 port map( G => n19, D => N196, Q => 
                           data2i_22_port);
   data2i_reg_21_inst : DLH_X1 port map( G => n19, D => N195, Q => 
                           data2i_21_port);
   data2i_reg_20_inst : DLH_X1 port map( G => n19, D => N194, Q => 
                           data2i_20_port);
   data2i_reg_19_inst : DLH_X1 port map( G => n19, D => N193, Q => 
                           data2i_19_port);
   data2i_reg_18_inst : DLH_X1 port map( G => n19, D => N192, Q => 
                           data2i_18_port);
   data2i_reg_17_inst : DLH_X1 port map( G => n19, D => N191, Q => 
                           data2i_17_port);
   data2i_reg_16_inst : DLH_X1 port map( G => n19, D => N190, Q => 
                           data2i_16_port);
   data2i_reg_15_inst : DLH_X1 port map( G => n19, D => N189, Q => 
                           data2i_15_port);
   data2i_reg_14_inst : DLH_X1 port map( G => n19, D => N188, Q => 
                           data2i_14_port);
   data2i_reg_13_inst : DLH_X1 port map( G => n19, D => N187, Q => 
                           data2i_13_port);
   data2i_reg_12_inst : DLH_X1 port map( G => n19, D => N186, Q => 
                           data2i_12_port);
   data2i_reg_11_inst : DLH_X1 port map( G => n19, D => N185, Q => 
                           data2i_11_port);
   data2i_reg_10_inst : DLH_X1 port map( G => n19, D => N184, Q => 
                           data2i_10_port);
   data2i_reg_9_inst : DLH_X1 port map( G => n19, D => N183, Q => data2i_9_port
                           );
   data2i_reg_8_inst : DLH_X1 port map( G => n20, D => N182, Q => data2i_8_port
                           );
   data2i_reg_7_inst : DLH_X1 port map( G => n20, D => N181, Q => data2i_7_port
                           );
   data2i_reg_6_inst : DLH_X1 port map( G => n20, D => N180, Q => data2i_6_port
                           );
   data2i_reg_5_inst : DLH_X1 port map( G => n20, D => N179, Q => data2i_5_port
                           );
   data2i_reg_4_inst : DLH_X1 port map( G => n20, D => N178, Q => data2i_4_port
                           );
   data2i_reg_3_inst : DLH_X1 port map( G => n20, D => N177, Q => data2i_3_port
                           );
   data2i_reg_2_inst : DLH_X1 port map( G => n20, D => N176, Q => data2i_2_port
                           );
   data2i_reg_1_inst : DLH_X1 port map( G => n20, D => N175, Q => data2i_1_port
                           );
   data2i_reg_0_inst : DLH_X1 port map( G => n20, D => N174, Q => data2i_0_port
                           );
   data1i_reg_31_inst : DLH_X1 port map( G => n20, D => DATA1(31), Q => 
                           data1i_31_port);
   data1i_reg_30_inst : DLH_X1 port map( G => n20, D => DATA1(30), Q => 
                           data1i_30_port);
   data1i_reg_29_inst : DLH_X1 port map( G => n20, D => DATA1(29), Q => 
                           data1i_29_port);
   data1i_reg_28_inst : DLH_X1 port map( G => n20, D => DATA1(28), Q => 
                           data1i_28_port);
   data1i_reg_27_inst : DLH_X1 port map( G => n20, D => DATA1(27), Q => 
                           data1i_27_port);
   data1i_reg_26_inst : DLH_X1 port map( G => n20, D => DATA1(26), Q => 
                           data1i_26_port);
   data1i_reg_25_inst : DLH_X1 port map( G => n20, D => DATA1(25), Q => 
                           data1i_25_port);
   data1i_reg_24_inst : DLH_X1 port map( G => n20, D => DATA1(24), Q => 
                           data1i_24_port);
   data1i_reg_23_inst : DLH_X1 port map( G => n20, D => DATA1(23), Q => 
                           data1i_23_port);
   data1i_reg_22_inst : DLH_X1 port map( G => n20, D => DATA1(22), Q => 
                           data1i_22_port);
   data1i_reg_21_inst : DLH_X1 port map( G => n20, D => DATA1(21), Q => 
                           data1i_21_port);
   data1i_reg_20_inst : DLH_X1 port map( G => n20, D => DATA1(20), Q => 
                           data1i_20_port);
   data1i_reg_19_inst : DLH_X1 port map( G => n20, D => DATA1(19), Q => 
                           data1i_19_port);
   data1i_reg_18_inst : DLH_X1 port map( G => n20, D => DATA1(18), Q => 
                           data1i_18_port);
   data1i_reg_17_inst : DLH_X1 port map( G => n20, D => DATA1(17), Q => 
                           data1i_17_port);
   data1i_reg_16_inst : DLH_X1 port map( G => n20, D => DATA1(16), Q => 
                           data1i_16_port);
   data1i_reg_15_inst : DLH_X1 port map( G => n20, D => DATA1(15), Q => 
                           data1i_15_port);
   data1i_reg_14_inst : DLH_X1 port map( G => n20, D => DATA1(14), Q => 
                           data1i_14_port);
   data1i_reg_13_inst : DLH_X1 port map( G => n21, D => DATA1(13), Q => 
                           data1i_13_port);
   data1i_reg_12_inst : DLH_X1 port map( G => n21, D => DATA1(12), Q => 
                           data1i_12_port);
   data1i_reg_11_inst : DLH_X1 port map( G => n21, D => DATA1(11), Q => 
                           data1i_11_port);
   data1i_reg_10_inst : DLH_X1 port map( G => n21, D => DATA1(10), Q => 
                           data1i_10_port);
   data1i_reg_9_inst : DLH_X1 port map( G => n21, D => DATA1(9), Q => 
                           data1i_9_port);
   data1i_reg_8_inst : DLH_X1 port map( G => n21, D => DATA1(8), Q => 
                           data1i_8_port);
   data1i_reg_7_inst : DLH_X1 port map( G => n21, D => DATA1(7), Q => 
                           data1i_7_port);
   data1i_reg_6_inst : DLH_X1 port map( G => n21, D => DATA1(6), Q => 
                           data1i_6_port);
   data1i_reg_5_inst : DLH_X1 port map( G => n21, D => DATA1(5), Q => 
                           data1i_5_port);
   data1i_reg_4_inst : DLH_X1 port map( G => n21, D => DATA1(4), Q => 
                           data1i_4_port);
   data1i_reg_3_inst : DLH_X1 port map( G => n21, D => DATA1(3), Q => 
                           data1i_3_port);
   data1i_reg_2_inst : DLH_X1 port map( G => n21, D => DATA1(2), Q => 
                           data1i_2_port);
   data1i_reg_1_inst : DLH_X1 port map( G => n21, D => DATA1(1), Q => 
                           data1i_1_port);
   data1i_reg_0_inst : DLH_X1 port map( G => n21, D => DATA1(0), Q => 
                           data1i_0_port);
   LOGIC_ARITH_i_reg : DLH_X1 port map( G => n15, D => n164_port, Q => 
                           LOGIC_ARITH_i);
   LEFT_RIGHT_i_reg : DLH_X1 port map( G => n15, D => n164_port, Q => 
                           LEFT_RIGHT_i);
   OUTPUT_alu_i_reg_0_inst : DLH_X1 port map( G => n16, D => N142, Q => 
                           OUTPUT_alu_i_0_port);
   OUT_ALU_reg_0_inst : DFF_X1 port map( D => OUTPUT_alu_i_0_port, CK => CLK, Q
                           => OUT_ALU(0), QN => n_1089);
   OUTPUT_alu_i_reg_1_inst : DLH_X1 port map( G => n16, D => N143, Q => 
                           OUTPUT_alu_i_1_port);
   OUT_ALU_reg_1_inst : DFF_X1 port map( D => OUTPUT_alu_i_1_port, CK => CLK, Q
                           => OUT_ALU(1), QN => n_1090);
   OUTPUT_alu_i_reg_2_inst : DLH_X1 port map( G => n16, D => N144, Q => 
                           OUTPUT_alu_i_2_port);
   OUT_ALU_reg_2_inst : DFF_X1 port map( D => OUTPUT_alu_i_2_port, CK => CLK, Q
                           => OUT_ALU(2), QN => n_1091);
   OUTPUT_alu_i_reg_3_inst : DLH_X1 port map( G => n16, D => N145, Q => 
                           OUTPUT_alu_i_3_port);
   OUT_ALU_reg_3_inst : DFF_X1 port map( D => OUTPUT_alu_i_3_port, CK => CLK, Q
                           => OUT_ALU(3), QN => n_1092);
   OUTPUT_alu_i_reg_4_inst : DLH_X1 port map( G => n16, D => N146, Q => 
                           OUTPUT_alu_i_4_port);
   OUT_ALU_reg_4_inst : DFF_X1 port map( D => OUTPUT_alu_i_4_port, CK => CLK, Q
                           => OUT_ALU(4), QN => n_1093);
   OUTPUT_alu_i_reg_5_inst : DLH_X1 port map( G => n16, D => N147, Q => 
                           OUTPUT_alu_i_5_port);
   OUT_ALU_reg_5_inst : DFF_X1 port map( D => OUTPUT_alu_i_5_port, CK => CLK, Q
                           => OUT_ALU(5), QN => n_1094);
   OUTPUT_alu_i_reg_6_inst : DLH_X1 port map( G => n16, D => N148, Q => 
                           OUTPUT_alu_i_6_port);
   OUT_ALU_reg_6_inst : DFF_X1 port map( D => OUTPUT_alu_i_6_port, CK => CLK, Q
                           => OUT_ALU(6), QN => n_1095);
   OUTPUT_alu_i_reg_7_inst : DLH_X1 port map( G => n16, D => N149, Q => 
                           OUTPUT_alu_i_7_port);
   OUT_ALU_reg_7_inst : DFF_X1 port map( D => OUTPUT_alu_i_7_port, CK => CLK, Q
                           => OUT_ALU(7), QN => n_1096);
   OUTPUT_alu_i_reg_8_inst : DLH_X1 port map( G => n16, D => N150, Q => 
                           OUTPUT_alu_i_8_port);
   OUT_ALU_reg_8_inst : DFF_X1 port map( D => OUTPUT_alu_i_8_port, CK => CLK, Q
                           => OUT_ALU(8), QN => n_1097);
   OUTPUT_alu_i_reg_9_inst : DLH_X1 port map( G => n16, D => N151, Q => 
                           OUTPUT_alu_i_9_port);
   OUT_ALU_reg_9_inst : DFF_X1 port map( D => OUTPUT_alu_i_9_port, CK => CLK, Q
                           => OUT_ALU(9), QN => n_1098);
   OUTPUT_alu_i_reg_10_inst : DLH_X1 port map( G => n16, D => N152, Q => 
                           OUTPUT_alu_i_10_port);
   OUT_ALU_reg_10_inst : DFF_X1 port map( D => OUTPUT_alu_i_10_port, CK => CLK,
                           Q => OUT_ALU(10), QN => n_1099);
   OUTPUT_alu_i_reg_11_inst : DLH_X1 port map( G => n17, D => N153, Q => 
                           OUTPUT_alu_i_11_port);
   OUT_ALU_reg_11_inst : DFF_X1 port map( D => OUTPUT_alu_i_11_port, CK => CLK,
                           Q => OUT_ALU(11), QN => n_1100);
   OUTPUT_alu_i_reg_12_inst : DLH_X1 port map( G => n17, D => N154, Q => 
                           OUTPUT_alu_i_12_port);
   OUT_ALU_reg_12_inst : DFF_X1 port map( D => OUTPUT_alu_i_12_port, CK => CLK,
                           Q => OUT_ALU(12), QN => n_1101);
   OUTPUT_alu_i_reg_13_inst : DLH_X1 port map( G => n17, D => N155, Q => 
                           OUTPUT_alu_i_13_port);
   OUT_ALU_reg_13_inst : DFF_X1 port map( D => OUTPUT_alu_i_13_port, CK => CLK,
                           Q => OUT_ALU(13), QN => n_1102);
   OUTPUT_alu_i_reg_14_inst : DLH_X1 port map( G => n17, D => N156, Q => 
                           OUTPUT_alu_i_14_port);
   OUT_ALU_reg_14_inst : DFF_X1 port map( D => OUTPUT_alu_i_14_port, CK => CLK,
                           Q => OUT_ALU(14), QN => n_1103);
   OUTPUT_alu_i_reg_15_inst : DLH_X1 port map( G => n17, D => N157, Q => 
                           OUTPUT_alu_i_15_port);
   OUT_ALU_reg_15_inst : DFF_X1 port map( D => OUTPUT_alu_i_15_port, CK => CLK,
                           Q => OUT_ALU(15), QN => n_1104);
   OUTPUT_alu_i_reg_16_inst : DLH_X1 port map( G => n17, D => N158, Q => 
                           OUTPUT_alu_i_16_port);
   OUT_ALU_reg_16_inst : DFF_X1 port map( D => OUTPUT_alu_i_16_port, CK => CLK,
                           Q => OUT_ALU(16), QN => n_1105);
   OUTPUT_alu_i_reg_17_inst : DLH_X1 port map( G => n17, D => N159, Q => 
                           OUTPUT_alu_i_17_port);
   OUT_ALU_reg_17_inst : DFF_X1 port map( D => OUTPUT_alu_i_17_port, CK => CLK,
                           Q => OUT_ALU(17), QN => n_1106);
   OUTPUT_alu_i_reg_18_inst : DLH_X1 port map( G => n17, D => N160, Q => 
                           OUTPUT_alu_i_18_port);
   OUT_ALU_reg_18_inst : DFF_X1 port map( D => OUTPUT_alu_i_18_port, CK => CLK,
                           Q => OUT_ALU(18), QN => n_1107);
   OUTPUT_alu_i_reg_19_inst : DLH_X1 port map( G => n17, D => N161, Q => 
                           OUTPUT_alu_i_19_port);
   OUT_ALU_reg_19_inst : DFF_X1 port map( D => OUTPUT_alu_i_19_port, CK => CLK,
                           Q => OUT_ALU(19), QN => n_1108);
   OUTPUT_alu_i_reg_20_inst : DLH_X1 port map( G => n17, D => N162, Q => 
                           OUTPUT_alu_i_20_port);
   OUT_ALU_reg_20_inst : DFF_X1 port map( D => OUTPUT_alu_i_20_port, CK => CLK,
                           Q => OUT_ALU(20), QN => n_1109);
   OUTPUT_alu_i_reg_21_inst : DLH_X1 port map( G => n17, D => N163, Q => 
                           OUTPUT_alu_i_21_port);
   OUT_ALU_reg_21_inst : DFF_X1 port map( D => OUTPUT_alu_i_21_port, CK => CLK,
                           Q => OUT_ALU(21), QN => n_1110);
   OUTPUT_alu_i_reg_22_inst : DLH_X1 port map( G => n18, D => N164, Q => 
                           OUTPUT_alu_i_22_port);
   OUT_ALU_reg_22_inst : DFF_X1 port map( D => OUTPUT_alu_i_22_port, CK => CLK,
                           Q => OUT_ALU(22), QN => n_1111);
   OUTPUT_alu_i_reg_23_inst : DLH_X1 port map( G => n18, D => N165, Q => 
                           OUTPUT_alu_i_23_port);
   OUT_ALU_reg_23_inst : DFF_X1 port map( D => OUTPUT_alu_i_23_port, CK => CLK,
                           Q => OUT_ALU(23), QN => n_1112);
   OUTPUT_alu_i_reg_24_inst : DLH_X1 port map( G => n18, D => N166, Q => 
                           OUTPUT_alu_i_24_port);
   OUT_ALU_reg_24_inst : DFF_X1 port map( D => OUTPUT_alu_i_24_port, CK => CLK,
                           Q => OUT_ALU(24), QN => n_1113);
   OUTPUT_alu_i_reg_25_inst : DLH_X1 port map( G => n18, D => N167, Q => 
                           OUTPUT_alu_i_25_port);
   OUT_ALU_reg_25_inst : DFF_X1 port map( D => OUTPUT_alu_i_25_port, CK => CLK,
                           Q => OUT_ALU(25), QN => n_1114);
   OUTPUT_alu_i_reg_26_inst : DLH_X1 port map( G => n18, D => N168, Q => 
                           OUTPUT_alu_i_26_port);
   OUT_ALU_reg_26_inst : DFF_X1 port map( D => OUTPUT_alu_i_26_port, CK => CLK,
                           Q => OUT_ALU(26), QN => n_1115);
   OUTPUT_alu_i_reg_27_inst : DLH_X1 port map( G => n18, D => N169, Q => 
                           OUTPUT_alu_i_27_port);
   OUT_ALU_reg_27_inst : DFF_X1 port map( D => OUTPUT_alu_i_27_port, CK => CLK,
                           Q => OUT_ALU(27), QN => n_1116);
   OUTPUT_alu_i_reg_28_inst : DLH_X1 port map( G => n18, D => N170, Q => 
                           OUTPUT_alu_i_28_port);
   OUT_ALU_reg_28_inst : DFF_X1 port map( D => OUTPUT_alu_i_28_port, CK => CLK,
                           Q => OUT_ALU(28), QN => n_1117);
   OUTPUT_alu_i_reg_29_inst : DLH_X1 port map( G => n18, D => N171, Q => 
                           OUTPUT_alu_i_29_port);
   OUT_ALU_reg_29_inst : DFF_X1 port map( D => OUTPUT_alu_i_29_port, CK => CLK,
                           Q => OUT_ALU(29), QN => n_1118);
   OUTPUT_alu_i_reg_30_inst : DLH_X1 port map( G => n18, D => N172, Q => 
                           OUTPUT_alu_i_30_port);
   OUT_ALU_reg_30_inst : DFF_X1 port map( D => OUTPUT_alu_i_30_port, CK => CLK,
                           Q => OUT_ALU(30), QN => n_1119);
   OUTPUT_alu_i_reg_31_inst : DLH_X1 port map( G => n18, D => N173, Q => 
                           OUTPUT_alu_i_31_port);
   OUT_ALU_reg_31_inst : DFF_X1 port map( D => OUTPUT_alu_i_31_port, CK => CLK,
                           Q => OUT_ALU(31), QN => n_1120);
   SHIFT_ROTATE_i <= '1';
   U221 : NAND3_X1 port map( A1 => n144_port, A2 => n143_port, A3 => n152_port,
                           ZN => n149_port);
   U222 : NAND3_X1 port map( A1 => n133, A2 => n168_port, A3 => FUNC(3), ZN => 
                           n143_port);
   U223 : NAND3_X1 port map( A1 => n147_port, A2 => n168_port, A3 => FUNC(3), 
                           ZN => n122);
   log : logic_N32 port map( FUNC(0) => FUNC(0), FUNC(1) => FUNC(1), FUNC(2) =>
                           FUNC(2), FUNC(3) => FUNC(3), FUNC(4) => FUNC(4), 
                           FUNC(5) => FUNC(5), DATA1(31) => DATA1(31), 
                           DATA1(30) => DATA1(30), DATA1(29) => DATA1(29), 
                           DATA1(28) => DATA1(28), DATA1(27) => DATA1(27), 
                           DATA1(26) => DATA1(26), DATA1(25) => DATA1(25), 
                           DATA1(24) => DATA1(24), DATA1(23) => DATA1(23), 
                           DATA1(22) => DATA1(22), DATA1(21) => DATA1(21), 
                           DATA1(20) => DATA1(20), DATA1(19) => DATA1(19), 
                           DATA1(18) => DATA1(18), DATA1(17) => DATA1(17), 
                           DATA1(16) => DATA1(16), DATA1(15) => DATA1(15), 
                           DATA1(14) => DATA1(14), DATA1(13) => DATA1(13), 
                           DATA1(12) => DATA1(12), DATA1(11) => DATA1(11), 
                           DATA1(10) => DATA1(10), DATA1(9) => DATA1(9), 
                           DATA1(8) => DATA1(8), DATA1(7) => DATA1(7), DATA1(6)
                           => DATA1(6), DATA1(5) => DATA1(5), DATA1(4) => 
                           DATA1(4), DATA1(3) => DATA1(3), DATA1(2) => DATA1(2)
                           , DATA1(1) => DATA1(1), DATA1(0) => DATA1(0), 
                           DATA2(31) => DATA2(31), DATA2(30) => DATA2(30), 
                           DATA2(29) => DATA2(29), DATA2(28) => DATA2(28), 
                           DATA2(27) => DATA2(27), DATA2(26) => DATA2(26), 
                           DATA2(25) => DATA2(25), DATA2(24) => DATA2(24), 
                           DATA2(23) => DATA2(23), DATA2(22) => DATA2(22), 
                           DATA2(21) => DATA2(21), DATA2(20) => DATA2(20), 
                           DATA2(19) => DATA2(19), DATA2(18) => DATA2(18), 
                           DATA2(17) => DATA2(17), DATA2(16) => DATA2(16), 
                           DATA2(15) => DATA2(15), DATA2(14) => DATA2(14), 
                           DATA2(13) => DATA2(13), DATA2(12) => DATA2(12), 
                           DATA2(11) => DATA2(11), DATA2(10) => DATA2(10), 
                           DATA2(9) => DATA2(9), DATA2(8) => DATA2(8), DATA2(7)
                           => DATA2(7), DATA2(6) => DATA2(6), DATA2(5) => 
                           DATA2(5), DATA2(4) => DATA2(4), DATA2(3) => n26, 
                           DATA2(2) => n24, DATA2(1) => DATA2(1), DATA2(0) => 
                           DATA2(0), OUT_ALU(31) => OUTPUT4_31_port, 
                           OUT_ALU(30) => OUTPUT4_30_port, OUT_ALU(29) => 
                           OUTPUT4_29_port, OUT_ALU(28) => OUTPUT4_28_port, 
                           OUT_ALU(27) => OUTPUT4_27_port, OUT_ALU(26) => 
                           OUTPUT4_26_port, OUT_ALU(25) => OUTPUT4_25_port, 
                           OUT_ALU(24) => OUTPUT4_24_port, OUT_ALU(23) => 
                           OUTPUT4_23_port, OUT_ALU(22) => OUTPUT4_22_port, 
                           OUT_ALU(21) => OUTPUT4_21_port, OUT_ALU(20) => 
                           OUTPUT4_20_port, OUT_ALU(19) => OUTPUT4_19_port, 
                           OUT_ALU(18) => OUTPUT4_18_port, OUT_ALU(17) => 
                           OUTPUT4_17_port, OUT_ALU(16) => OUTPUT4_16_port, 
                           OUT_ALU(15) => OUTPUT4_15_port, OUT_ALU(14) => 
                           OUTPUT4_14_port, OUT_ALU(13) => OUTPUT4_13_port, 
                           OUT_ALU(12) => OUTPUT4_12_port, OUT_ALU(11) => 
                           OUTPUT4_11_port, OUT_ALU(10) => OUTPUT4_10_port, 
                           OUT_ALU(9) => OUTPUT4_9_port, OUT_ALU(8) => 
                           OUTPUT4_8_port, OUT_ALU(7) => OUTPUT4_7_port, 
                           OUT_ALU(6) => OUTPUT4_6_port, OUT_ALU(5) => 
                           OUTPUT4_5_port, OUT_ALU(4) => OUTPUT4_4_port, 
                           OUT_ALU(3) => OUTPUT4_3_port, OUT_ALU(2) => 
                           OUTPUT4_2_port, OUT_ALU(1) => OUTPUT4_1_port, 
                           OUT_ALU(0) => OUTPUT4_0_port);
   comp : comparator port map( DATA1(31) => OUTPUT2_31_port, DATA1(30) => 
                           OUTPUT2_30_port, DATA1(29) => OUTPUT2_29_port, 
                           DATA1(28) => OUTPUT2_28_port, DATA1(27) => 
                           OUTPUT2_27_port, DATA1(26) => OUTPUT2_26_port, 
                           DATA1(25) => OUTPUT2_25_port, DATA1(24) => 
                           OUTPUT2_24_port, DATA1(23) => OUTPUT2_23_port, 
                           DATA1(22) => OUTPUT2_22_port, DATA1(21) => 
                           OUTPUT2_21_port, DATA1(20) => OUTPUT2_20_port, 
                           DATA1(19) => OUTPUT2_19_port, DATA1(18) => 
                           OUTPUT2_18_port, DATA1(17) => OUTPUT2_17_port, 
                           DATA1(16) => OUTPUT2_16_port, DATA1(15) => 
                           OUTPUT2_15_port, DATA1(14) => OUTPUT2_14_port, 
                           DATA1(13) => OUTPUT2_13_port, DATA1(12) => 
                           OUTPUT2_12_port, DATA1(11) => OUTPUT2_11_port, 
                           DATA1(10) => OUTPUT2_10_port, DATA1(9) => 
                           OUTPUT2_9_port, DATA1(8) => OUTPUT2_8_port, DATA1(7)
                           => OUTPUT2_7_port, DATA1(6) => OUTPUT2_6_port, 
                           DATA1(5) => OUTPUT2_5_port, DATA1(4) => 
                           OUTPUT2_4_port, DATA1(3) => OUTPUT2_3_port, DATA1(2)
                           => OUTPUT2_2_port, DATA1(1) => OUTPUT2_1_port, 
                           DATA1(0) => OUTPUT2_0_port, DATA2i => Cout_i, 
                           tipo(0) => FUNC(0), tipo(1) => FUNC(1), tipo(2) => 
                           FUNC(2), tipo(3) => FUNC(3), tipo(4) => FUNC(4), 
                           tipo(5) => FUNC(5), OUTALU(31) => n_1121, OUTALU(30)
                           => n_1122, OUTALU(29) => n_1123, OUTALU(28) => 
                           n_1124, OUTALU(27) => n_1125, OUTALU(26) => n_1126, 
                           OUTALU(25) => n_1127, OUTALU(24) => n_1128, 
                           OUTALU(23) => n_1129, OUTALU(22) => n_1130, 
                           OUTALU(21) => n_1131, OUTALU(20) => n_1132, 
                           OUTALU(19) => n_1133, OUTALU(18) => n_1134, 
                           OUTALU(17) => n_1135, OUTALU(16) => n_1136, 
                           OUTALU(15) => n_1137, OUTALU(14) => n_1138, 
                           OUTALU(13) => n_1139, OUTALU(12) => n_1140, 
                           OUTALU(11) => n_1141, OUTALU(10) => n_1142, 
                           OUTALU(9) => n_1143, OUTALU(8) => n_1144, OUTALU(7) 
                           => n_1145, OUTALU(6) => n_1146, OUTALU(5) => n_1147,
                           OUTALU(4) => n_1148, OUTALU(3) => n_1149, OUTALU(2) 
                           => n_1150, OUTALU(1) => n_1151, OUTALU(0) => 
                           OUTPUT3_0_port);
   shifter : SHIFTER_GENERIC_N32 port map( A(31) => DATA1(31), A(30) => 
                           DATA1(30), A(29) => DATA1(29), A(28) => DATA1(28), 
                           A(27) => DATA1(27), A(26) => DATA1(26), A(25) => 
                           DATA1(25), A(24) => DATA1(24), A(23) => DATA1(23), 
                           A(22) => DATA1(22), A(21) => DATA1(21), A(20) => 
                           DATA1(20), A(19) => DATA1(19), A(18) => DATA1(18), 
                           A(17) => DATA1(17), A(16) => DATA1(16), A(15) => 
                           DATA1(15), A(14) => DATA1(14), A(13) => DATA1(13), 
                           A(12) => DATA1(12), A(11) => DATA1(11), A(10) => 
                           DATA1(10), A(9) => DATA1(9), A(8) => DATA1(8), A(7) 
                           => DATA1(7), A(6) => DATA1(6), A(5) => DATA1(5), 
                           A(4) => DATA1(4), A(3) => DATA1(3), A(2) => DATA1(2)
                           , A(1) => DATA1(1), A(0) => DATA1(0), B(4) => 
                           DATA2(4), B(3) => n26, B(2) => n24, B(1) => DATA2(1)
                           , B(0) => DATA2(0), LOGIC_ARITH => LOGIC_ARITH_i, 
                           LEFT_RIGHT => LEFT_RIGHT_i, SHIFT_ROTATE => 
                           SHIFT_ROTATE_i, OUTPUT(31) => OUTPUT1_31_port, 
                           OUTPUT(30) => OUTPUT1_30_port, OUTPUT(29) => 
                           OUTPUT1_29_port, OUTPUT(28) => OUTPUT1_28_port, 
                           OUTPUT(27) => OUTPUT1_27_port, OUTPUT(26) => 
                           OUTPUT1_26_port, OUTPUT(25) => OUTPUT1_25_port, 
                           OUTPUT(24) => OUTPUT1_24_port, OUTPUT(23) => 
                           OUTPUT1_23_port, OUTPUT(22) => OUTPUT1_22_port, 
                           OUTPUT(21) => OUTPUT1_21_port, OUTPUT(20) => 
                           OUTPUT1_20_port, OUTPUT(19) => OUTPUT1_19_port, 
                           OUTPUT(18) => OUTPUT1_18_port, OUTPUT(17) => 
                           OUTPUT1_17_port, OUTPUT(16) => OUTPUT1_16_port, 
                           OUTPUT(15) => OUTPUT1_15_port, OUTPUT(14) => 
                           OUTPUT1_14_port, OUTPUT(13) => OUTPUT1_13_port, 
                           OUTPUT(12) => OUTPUT1_12_port, OUTPUT(11) => 
                           OUTPUT1_11_port, OUTPUT(10) => OUTPUT1_10_port, 
                           OUTPUT(9) => OUTPUT1_9_port, OUTPUT(8) => 
                           OUTPUT1_8_port, OUTPUT(7) => OUTPUT1_7_port, 
                           OUTPUT(6) => OUTPUT1_6_port, OUTPUT(5) => 
                           OUTPUT1_5_port, OUTPUT(4) => OUTPUT1_4_port, 
                           OUTPUT(3) => OUTPUT1_3_port, OUTPUT(2) => 
                           OUTPUT1_2_port, OUTPUT(1) => OUTPUT1_1_port, 
                           OUTPUT(0) => OUTPUT1_0_port);
   adder : P4_ADDER_NBIT32 port map( A(31) => data1i_31_port, A(30) => 
                           data1i_30_port, A(29) => data1i_29_port, A(28) => 
                           data1i_28_port, A(27) => data1i_27_port, A(26) => 
                           data1i_26_port, A(25) => data1i_25_port, A(24) => 
                           data1i_24_port, A(23) => data1i_23_port, A(22) => 
                           data1i_22_port, A(21) => data1i_21_port, A(20) => 
                           data1i_20_port, A(19) => data1i_19_port, A(18) => 
                           data1i_18_port, A(17) => data1i_17_port, A(16) => 
                           data1i_16_port, A(15) => data1i_15_port, A(14) => 
                           data1i_14_port, A(13) => data1i_13_port, A(12) => 
                           data1i_12_port, A(11) => data1i_11_port, A(10) => 
                           data1i_10_port, A(9) => data1i_9_port, A(8) => 
                           data1i_8_port, A(7) => data1i_7_port, A(6) => 
                           data1i_6_port, A(5) => data1i_5_port, A(4) => 
                           data1i_4_port, A(3) => data1i_3_port, A(2) => 
                           data1i_2_port, A(1) => data1i_1_port, A(0) => 
                           data1i_0_port, B(31) => data2i_31_port, B(30) => 
                           data2i_30_port, B(29) => data2i_29_port, B(28) => 
                           data2i_28_port, B(27) => data2i_27_port, B(26) => 
                           data2i_26_port, B(25) => data2i_25_port, B(24) => 
                           data2i_24_port, B(23) => data2i_23_port, B(22) => 
                           data2i_22_port, B(21) => data2i_21_port, B(20) => 
                           data2i_20_port, B(19) => data2i_19_port, B(18) => 
                           data2i_18_port, B(17) => data2i_17_port, B(16) => 
                           data2i_16_port, B(15) => data2i_15_port, B(14) => 
                           data2i_14_port, B(13) => data2i_13_port, B(12) => 
                           data2i_12_port, B(11) => data2i_11_port, B(10) => 
                           data2i_10_port, B(9) => data2i_9_port, B(8) => 
                           data2i_8_port, B(7) => data2i_7_port, B(6) => 
                           data2i_6_port, B(5) => data2i_5_port, B(4) => 
                           data2i_4_port, B(3) => data2i_3_port, B(2) => 
                           data2i_2_port, B(1) => data2i_1_port, B(0) => 
                           data2i_0_port, Cin => Cin_i, S(31) => 
                           OUTPUT2_31_port, S(30) => OUTPUT2_30_port, S(29) => 
                           OUTPUT2_29_port, S(28) => OUTPUT2_28_port, S(27) => 
                           OUTPUT2_27_port, S(26) => OUTPUT2_26_port, S(25) => 
                           OUTPUT2_25_port, S(24) => OUTPUT2_24_port, S(23) => 
                           OUTPUT2_23_port, S(22) => OUTPUT2_22_port, S(21) => 
                           OUTPUT2_21_port, S(20) => OUTPUT2_20_port, S(19) => 
                           OUTPUT2_19_port, S(18) => OUTPUT2_18_port, S(17) => 
                           OUTPUT2_17_port, S(16) => OUTPUT2_16_port, S(15) => 
                           OUTPUT2_15_port, S(14) => OUTPUT2_14_port, S(13) => 
                           OUTPUT2_13_port, S(12) => OUTPUT2_12_port, S(11) => 
                           OUTPUT2_11_port, S(10) => OUTPUT2_10_port, S(9) => 
                           OUTPUT2_9_port, S(8) => OUTPUT2_8_port, S(7) => 
                           OUTPUT2_7_port, S(6) => OUTPUT2_6_port, S(5) => 
                           OUTPUT2_5_port, S(4) => OUTPUT2_4_port, S(3) => 
                           OUTPUT2_3_port, S(2) => OUTPUT2_2_port, S(1) => 
                           OUTPUT2_1_port, S(0) => OUTPUT2_0_port, Cout => 
                           Cout_i);
   U4 : BUF_X1 port map( A => N139, Z => n20);
   U5 : BUF_X1 port map( A => n53, Z => n8);
   U6 : BUF_X1 port map( A => n53, Z => n9);
   U7 : INV_X1 port map( A => n1, ZN => n11);
   U8 : INV_X1 port map( A => n1, ZN => n12);
   U9 : BUF_X1 port map( A => N139, Z => n19);
   U10 : BUF_X1 port map( A => n162_port, Z => n2);
   U11 : BUF_X1 port map( A => n162_port, Z => n3);
   U12 : BUF_X1 port map( A => n162_port, Z => n4);
   U13 : BUF_X1 port map( A => n53, Z => n10);
   U14 : BUF_X1 port map( A => N139, Z => n21);
   U15 : BUF_X1 port map( A => N141, Z => n17);
   U16 : BUF_X1 port map( A => N141, Z => n16);
   U17 : BUF_X1 port map( A => N141, Z => n18);
   U18 : AOI21_X1 port map( B1 => n152_port, B2 => n120, A => n171_port, ZN => 
                           n134);
   U19 : BUF_X1 port map( A => n54, Z => n5);
   U20 : BUF_X1 port map( A => n54, Z => n6);
   U21 : BUF_X1 port map( A => n54, Z => n7);
   U22 : OR3_X1 port map( A1 => n134, A2 => n135, A3 => n55, ZN => n1);
   U23 : INV_X1 port map( A => n50, ZN => n162_port);
   U24 : NAND2_X1 port map( A1 => n132, A2 => n123, ZN => n130);
   U25 : NAND2_X1 port map( A1 => n124, A2 => n171_port, ZN => n140);
   U26 : OR3_X1 port map( A1 => n134, A2 => n135, A3 => n50, ZN => n53);
   U27 : OR2_X1 port map( A1 => n10, A2 => n55, ZN => N139);
   U28 : OR3_X1 port map( A1 => n19, A2 => n15, A3 => n7, ZN => N141);
   U29 : INV_X1 port map( A => n142_port, ZN => n167_port);
   U30 : NAND2_X1 port map( A1 => n51, A2 => n52, ZN => N173);
   U31 : NAND2_X1 port map( A1 => OUTPUT1_31_port, A2 => n13, ZN => n51);
   U32 : AOI22_X1 port map( A1 => OUTPUT2_31_port, A2 => n8, B1 => 
                           OUTPUT4_31_port, B2 => n5, ZN => n52);
   U33 : NAND2_X1 port map( A1 => n56, A2 => n57, ZN => N172);
   U34 : NAND2_X1 port map( A1 => OUTPUT1_30_port, A2 => n15, ZN => n56);
   U35 : AOI22_X1 port map( A1 => OUTPUT2_30_port, A2 => n8, B1 => 
                           OUTPUT4_30_port, B2 => n5, ZN => n57);
   U36 : NAND2_X1 port map( A1 => n58, A2 => n59, ZN => N171);
   U37 : NAND2_X1 port map( A1 => OUTPUT1_29_port, A2 => n15, ZN => n58);
   U38 : AOI22_X1 port map( A1 => OUTPUT2_29_port, A2 => n8, B1 => 
                           OUTPUT4_29_port, B2 => n5, ZN => n59);
   U39 : NAND2_X1 port map( A1 => n60, A2 => n61, ZN => N170);
   U40 : NAND2_X1 port map( A1 => OUTPUT1_28_port, A2 => n15, ZN => n60);
   U41 : AOI22_X1 port map( A1 => OUTPUT2_28_port, A2 => n8, B1 => 
                           OUTPUT4_28_port, B2 => n5, ZN => n61);
   U42 : NAND2_X1 port map( A1 => n62, A2 => n63, ZN => N169);
   U43 : NAND2_X1 port map( A1 => OUTPUT1_27_port, A2 => n15, ZN => n62);
   U44 : AOI22_X1 port map( A1 => OUTPUT2_27_port, A2 => n8, B1 => 
                           OUTPUT4_27_port, B2 => n5, ZN => n63);
   U45 : NAND2_X1 port map( A1 => n64, A2 => n65, ZN => N168);
   U46 : NAND2_X1 port map( A1 => OUTPUT1_26_port, A2 => n15, ZN => n64);
   U47 : AOI22_X1 port map( A1 => OUTPUT2_26_port, A2 => n8, B1 => 
                           OUTPUT4_26_port, B2 => n5, ZN => n65);
   U48 : NAND2_X1 port map( A1 => n66, A2 => n67, ZN => N167);
   U49 : NAND2_X1 port map( A1 => OUTPUT1_25_port, A2 => n15, ZN => n66);
   U50 : AOI22_X1 port map( A1 => OUTPUT2_25_port, A2 => n8, B1 => 
                           OUTPUT4_25_port, B2 => n5, ZN => n67);
   U51 : NAND2_X1 port map( A1 => n68, A2 => n69, ZN => N166);
   U52 : NAND2_X1 port map( A1 => OUTPUT1_24_port, A2 => n15, ZN => n68);
   U53 : AOI22_X1 port map( A1 => OUTPUT2_24_port, A2 => n8, B1 => 
                           OUTPUT4_24_port, B2 => n5, ZN => n69);
   U54 : NAND2_X1 port map( A1 => n70, A2 => n71, ZN => N165);
   U55 : NAND2_X1 port map( A1 => OUTPUT1_23_port, A2 => n14, ZN => n70);
   U56 : AOI22_X1 port map( A1 => OUTPUT2_23_port, A2 => n8, B1 => 
                           OUTPUT4_23_port, B2 => n5, ZN => n71);
   U57 : NAND2_X1 port map( A1 => n72, A2 => n73, ZN => N164);
   U58 : NAND2_X1 port map( A1 => OUTPUT1_22_port, A2 => n14, ZN => n72);
   U59 : AOI22_X1 port map( A1 => OUTPUT2_22_port, A2 => n8, B1 => 
                           OUTPUT4_22_port, B2 => n5, ZN => n73);
   U60 : NAND2_X1 port map( A1 => n74, A2 => n75, ZN => N163);
   U61 : NAND2_X1 port map( A1 => OUTPUT1_21_port, A2 => n14, ZN => n74);
   U62 : AOI22_X1 port map( A1 => OUTPUT2_21_port, A2 => n8, B1 => 
                           OUTPUT4_21_port, B2 => n5, ZN => n75);
   U63 : NAND2_X1 port map( A1 => n76, A2 => n77, ZN => N162);
   U64 : NAND2_X1 port map( A1 => OUTPUT1_20_port, A2 => n14, ZN => n76);
   U65 : AOI22_X1 port map( A1 => OUTPUT2_20_port, A2 => n8, B1 => 
                           OUTPUT4_20_port, B2 => n5, ZN => n77);
   U66 : NAND2_X1 port map( A1 => n78, A2 => n79, ZN => N161);
   U67 : NAND2_X1 port map( A1 => OUTPUT1_19_port, A2 => n14, ZN => n78);
   U68 : AOI22_X1 port map( A1 => OUTPUT2_19_port, A2 => n9, B1 => 
                           OUTPUT4_19_port, B2 => n6, ZN => n79);
   U69 : NAND2_X1 port map( A1 => n80, A2 => n81, ZN => N160);
   U70 : NAND2_X1 port map( A1 => OUTPUT1_18_port, A2 => n14, ZN => n80);
   U71 : AOI22_X1 port map( A1 => OUTPUT2_18_port, A2 => n9, B1 => 
                           OUTPUT4_18_port, B2 => n6, ZN => n81);
   U72 : NAND2_X1 port map( A1 => n82, A2 => n83, ZN => N159);
   U73 : NAND2_X1 port map( A1 => OUTPUT1_17_port, A2 => n14, ZN => n82);
   U74 : AOI22_X1 port map( A1 => OUTPUT2_17_port, A2 => n9, B1 => 
                           OUTPUT4_17_port, B2 => n6, ZN => n83);
   U75 : NAND2_X1 port map( A1 => n84, A2 => n85, ZN => N158);
   U76 : NAND2_X1 port map( A1 => OUTPUT1_16_port, A2 => n14, ZN => n84);
   U77 : AOI22_X1 port map( A1 => OUTPUT2_16_port, A2 => n9, B1 => 
                           OUTPUT4_16_port, B2 => n6, ZN => n85);
   U78 : NAND2_X1 port map( A1 => n86, A2 => n87, ZN => N157);
   U79 : NAND2_X1 port map( A1 => OUTPUT1_15_port, A2 => n14, ZN => n86);
   U80 : AOI22_X1 port map( A1 => OUTPUT2_15_port, A2 => n9, B1 => 
                           OUTPUT4_15_port, B2 => n6, ZN => n87);
   U81 : NAND2_X1 port map( A1 => n88, A2 => n89, ZN => N156);
   U82 : NAND2_X1 port map( A1 => OUTPUT1_14_port, A2 => n14, ZN => n88);
   U83 : AOI22_X1 port map( A1 => OUTPUT2_14_port, A2 => n9, B1 => 
                           OUTPUT4_14_port, B2 => n6, ZN => n89);
   U84 : NAND2_X1 port map( A1 => n90, A2 => n91, ZN => N155);
   U85 : NAND2_X1 port map( A1 => OUTPUT1_13_port, A2 => n14, ZN => n90);
   U86 : AOI22_X1 port map( A1 => OUTPUT2_13_port, A2 => n9, B1 => 
                           OUTPUT4_13_port, B2 => n6, ZN => n91);
   U87 : NAND2_X1 port map( A1 => n92, A2 => n93, ZN => N154);
   U88 : NAND2_X1 port map( A1 => OUTPUT1_12_port, A2 => n13, ZN => n92);
   U89 : AOI22_X1 port map( A1 => OUTPUT2_12_port, A2 => n9, B1 => 
                           OUTPUT4_12_port, B2 => n6, ZN => n93);
   U90 : NAND2_X1 port map( A1 => n94, A2 => n95, ZN => N153);
   U91 : NAND2_X1 port map( A1 => OUTPUT1_11_port, A2 => n13, ZN => n94);
   U92 : AOI22_X1 port map( A1 => OUTPUT2_11_port, A2 => n9, B1 => 
                           OUTPUT4_11_port, B2 => n6, ZN => n95);
   U93 : NAND2_X1 port map( A1 => n96, A2 => n97, ZN => N152);
   U94 : NAND2_X1 port map( A1 => OUTPUT1_10_port, A2 => n13, ZN => n96);
   U95 : AOI22_X1 port map( A1 => OUTPUT2_10_port, A2 => n9, B1 => 
                           OUTPUT4_10_port, B2 => n6, ZN => n97);
   U96 : NAND2_X1 port map( A1 => n98, A2 => n99, ZN => N151);
   U97 : NAND2_X1 port map( A1 => OUTPUT1_9_port, A2 => n13, ZN => n98);
   U98 : AOI22_X1 port map( A1 => OUTPUT2_9_port, A2 => n9, B1 => 
                           OUTPUT4_9_port, B2 => n6, ZN => n99);
   U99 : NAND2_X1 port map( A1 => n100, A2 => n101, ZN => N150);
   U100 : NAND2_X1 port map( A1 => OUTPUT1_8_port, A2 => n13, ZN => n100);
   U101 : AOI22_X1 port map( A1 => OUTPUT2_8_port, A2 => n9, B1 => 
                           OUTPUT4_8_port, B2 => n6, ZN => n101);
   U102 : NAND2_X1 port map( A1 => n102, A2 => n103, ZN => N149);
   U103 : NAND2_X1 port map( A1 => OUTPUT1_7_port, A2 => n13, ZN => n102);
   U104 : AOI22_X1 port map( A1 => OUTPUT2_7_port, A2 => n10, B1 => 
                           OUTPUT4_7_port, B2 => n7, ZN => n103);
   U105 : NAND2_X1 port map( A1 => n104, A2 => n105, ZN => N148);
   U106 : NAND2_X1 port map( A1 => OUTPUT1_6_port, A2 => n13, ZN => n104);
   U107 : AOI22_X1 port map( A1 => OUTPUT2_6_port, A2 => n10, B1 => 
                           OUTPUT4_6_port, B2 => n7, ZN => n105);
   U108 : NAND2_X1 port map( A1 => n106, A2 => n107, ZN => N147);
   U109 : NAND2_X1 port map( A1 => OUTPUT1_5_port, A2 => n14, ZN => n106);
   U110 : AOI22_X1 port map( A1 => OUTPUT2_5_port, A2 => n10, B1 => 
                           OUTPUT4_5_port, B2 => n7, ZN => n107);
   U111 : NAND2_X1 port map( A1 => n108, A2 => n109, ZN => N146);
   U112 : NAND2_X1 port map( A1 => OUTPUT1_4_port, A2 => n13, ZN => n108);
   U113 : AOI22_X1 port map( A1 => OUTPUT2_4_port, A2 => n10, B1 => 
                           OUTPUT4_4_port, B2 => n7, ZN => n109);
   U114 : INV_X1 port map( A => n48, ZN => n164_port);
   U115 : INV_X1 port map( A => n27, ZN => n26);
   U116 : OAI221_X1 port map( B1 => n173_port, B2 => n118, C1 => n119, C2 => 
                           n120, A => n165_port, ZN => n54);
   U117 : INV_X1 port map( A => n121, ZN => n165_port);
   U118 : OAI22_X1 port map( A1 => n122, A2 => n170_port, B1 => n123, B2 => 
                           n124, ZN => n121);
   U119 : INV_X1 port map( A => n125, ZN => n170_port);
   U120 : OAI221_X1 port map( B1 => n127, B2 => n118, C1 => n119, C2 => n136, A
                           => n137, ZN => n55);
   U121 : AOI221_X1 port map( B1 => n138, B2 => n125, C1 => n139_port, C2 => 
                           n140, A => n141_port, ZN => n137);
   U122 : NAND2_X1 port map( A1 => n143_port, A2 => n144_port, ZN => n139_port)
                           ;
   U123 : OAI211_X1 port map( C1 => n142_port, C2 => n161_port, A => n118, B =>
                           n126, ZN => n138);
   U124 : OAI221_X1 port map( B1 => n124, B2 => n120, C1 => n127, C2 => n132, A
                           => n148_port, ZN => n50);
   U125 : AOI222_X1 port map( A1 => n163_port, A2 => n140, B1 => n174_port, B2 
                           => n149_port, C1 => n150_port, C2 => n151_port, ZN 
                           => n148_port);
   U126 : INV_X1 port map( A => n136, ZN => n163_port);
   U127 : NOR2_X1 port map( A1 => n168_port, A2 => n169_port, ZN => n153_port);
   U128 : BUF_X1 port map( A => N206, Z => n15);
   U129 : AOI21_X1 port map( B1 => n122, B2 => n152_port, A => n127, ZN => n135
                           );
   U130 : BUF_X1 port map( A => N206, Z => n14);
   U131 : BUF_X1 port map( A => N206, Z => n13);
   U132 : NOR3_X1 port map( A1 => n166_port, A2 => n124, A3 => n142_port, ZN =>
                           n141_port);
   U133 : OAI22_X1 port map( A1 => DATA2(1), A2 => n11, B1 => n2, B2 => n23, ZN
                           => N175);
   U134 : OAI22_X1 port map( A1 => n24, A2 => n11, B1 => n2, B2 => n25, ZN => 
                           N176);
   U135 : OAI22_X1 port map( A1 => DATA2(0), A2 => n11, B1 => n2, B2 => n22, ZN
                           => N174);
   U136 : OAI22_X1 port map( A1 => DATA2(24), A2 => n11, B1 => n4, B2 => n36, 
                           ZN => N198);
   U137 : INV_X1 port map( A => DATA2(24), ZN => n36);
   U138 : OAI22_X1 port map( A1 => DATA2(25), A2 => n12, B1 => n4, B2 => n35, 
                           ZN => N199);
   U139 : INV_X1 port map( A => DATA2(25), ZN => n35);
   U140 : OAI22_X1 port map( A1 => DATA2(26), A2 => n11, B1 => n4, B2 => n34, 
                           ZN => N200);
   U141 : INV_X1 port map( A => DATA2(26), ZN => n34);
   U142 : OAI22_X1 port map( A1 => DATA2(27), A2 => n12, B1 => n4, B2 => n33, 
                           ZN => N201);
   U143 : INV_X1 port map( A => DATA2(27), ZN => n33);
   U144 : OAI22_X1 port map( A1 => DATA2(28), A2 => n11, B1 => n4, B2 => n32, 
                           ZN => N202);
   U145 : INV_X1 port map( A => DATA2(28), ZN => n32);
   U146 : OAI22_X1 port map( A1 => DATA2(29), A2 => n12, B1 => n4, B2 => n31, 
                           ZN => N203);
   U147 : INV_X1 port map( A => DATA2(29), ZN => n31);
   U148 : OAI22_X1 port map( A1 => DATA2(30), A2 => n11, B1 => n4, B2 => n30, 
                           ZN => N204);
   U149 : INV_X1 port map( A => DATA2(30), ZN => n30);
   U150 : OAI22_X1 port map( A1 => DATA2(31), A2 => n12, B1 => n4, B2 => n29, 
                           ZN => N205);
   U151 : INV_X1 port map( A => DATA2(31), ZN => n29);
   U152 : OAI22_X1 port map( A1 => n26, A2 => n11, B1 => n2, B2 => n27, ZN => 
                           N177);
   U153 : OAI22_X1 port map( A1 => DATA2(4), A2 => n11, B1 => n2, B2 => n28, ZN
                           => N178);
   U154 : OAI22_X1 port map( A1 => DATA2(5), A2 => n11, B1 => n2, B2 => 
                           n160_port, ZN => N179);
   U155 : INV_X1 port map( A => DATA2(5), ZN => n160_port);
   U156 : OAI22_X1 port map( A1 => DATA2(6), A2 => n11, B1 => n2, B2 => 
                           n159_port, ZN => N180);
   U157 : INV_X1 port map( A => DATA2(6), ZN => n159_port);
   U158 : OAI22_X1 port map( A1 => DATA2(7), A2 => n11, B1 => n2, B2 => 
                           n158_port, ZN => N181);
   U159 : INV_X1 port map( A => DATA2(7), ZN => n158_port);
   U160 : OAI22_X1 port map( A1 => DATA2(8), A2 => n11, B1 => n2, B2 => 
                           n157_port, ZN => N182);
   U161 : INV_X1 port map( A => DATA2(8), ZN => n157_port);
   U162 : OAI22_X1 port map( A1 => DATA2(9), A2 => n11, B1 => n2, B2 => 
                           n156_port, ZN => N183);
   U163 : INV_X1 port map( A => DATA2(9), ZN => n156_port);
   U164 : OAI22_X1 port map( A1 => DATA2(10), A2 => n11, B1 => n2, B2 => 
                           n155_port, ZN => N184);
   U165 : INV_X1 port map( A => DATA2(10), ZN => n155_port);
   U166 : OAI22_X1 port map( A1 => DATA2(11), A2 => n11, B1 => n2, B2 => 
                           n154_port, ZN => N185);
   U167 : INV_X1 port map( A => DATA2(11), ZN => n154_port);
   U168 : OAI22_X1 port map( A1 => DATA2(12), A2 => n12, B1 => n3, B2 => n49, 
                           ZN => N186);
   U169 : INV_X1 port map( A => DATA2(12), ZN => n49);
   U170 : OAI22_X1 port map( A1 => DATA2(13), A2 => n12, B1 => n3, B2 => n47, 
                           ZN => N187);
   U171 : INV_X1 port map( A => DATA2(13), ZN => n47);
   U172 : OAI22_X1 port map( A1 => DATA2(14), A2 => n12, B1 => n3, B2 => n46, 
                           ZN => N188);
   U173 : INV_X1 port map( A => DATA2(14), ZN => n46);
   U174 : OAI22_X1 port map( A1 => DATA2(15), A2 => n12, B1 => n3, B2 => n45, 
                           ZN => N189);
   U175 : INV_X1 port map( A => DATA2(15), ZN => n45);
   U176 : OAI22_X1 port map( A1 => DATA2(16), A2 => n12, B1 => n3, B2 => n44, 
                           ZN => N190);
   U177 : INV_X1 port map( A => DATA2(16), ZN => n44);
   U178 : OAI22_X1 port map( A1 => DATA2(17), A2 => n12, B1 => n3, B2 => n43, 
                           ZN => N191);
   U179 : INV_X1 port map( A => DATA2(17), ZN => n43);
   U180 : OAI22_X1 port map( A1 => DATA2(18), A2 => n12, B1 => n3, B2 => n42, 
                           ZN => N192);
   U181 : INV_X1 port map( A => DATA2(18), ZN => n42);
   U182 : OAI22_X1 port map( A1 => DATA2(19), A2 => n12, B1 => n3, B2 => n41, 
                           ZN => N193);
   U183 : INV_X1 port map( A => DATA2(19), ZN => n41);
   U184 : OAI22_X1 port map( A1 => DATA2(20), A2 => n12, B1 => n3, B2 => n40, 
                           ZN => N194);
   U185 : INV_X1 port map( A => DATA2(20), ZN => n40);
   U186 : OAI22_X1 port map( A1 => DATA2(21), A2 => n12, B1 => n3, B2 => n39, 
                           ZN => N195);
   U187 : INV_X1 port map( A => DATA2(21), ZN => n39);
   U188 : OAI22_X1 port map( A1 => DATA2(22), A2 => n12, B1 => n3, B2 => n38, 
                           ZN => N196);
   U189 : INV_X1 port map( A => DATA2(22), ZN => n38);
   U190 : OAI22_X1 port map( A1 => DATA2(23), A2 => n12, B1 => n3, B2 => n37, 
                           ZN => N197);
   U191 : INV_X1 port map( A => DATA2(23), ZN => n37);
   U192 : NAND2_X1 port map( A1 => n146_port, A2 => n133, ZN => n152_port);
   U193 : AND2_X1 port map( A1 => n127, A2 => n173_port, ZN => n124);
   U194 : NAND4_X1 port map( A1 => n122, A2 => n152_port, A3 => n126, A4 => 
                           n132, ZN => n151_port);
   U195 : NAND2_X1 port map( A1 => n153_port, A2 => n147_port, ZN => n120);
   U196 : NAND2_X1 port map( A1 => n168_port, A2 => n169_port, ZN => n142_port)
                           ;
   U197 : NAND2_X1 port map( A1 => n146_port, A2 => n147_port, ZN => n118);
   U198 : NAND2_X1 port map( A1 => n147_port, A2 => n167_port, ZN => n132);
   U199 : NAND2_X1 port map( A1 => n153_port, A2 => n133, ZN => n126);
   U200 : INV_X1 port map( A => n129, ZN => n171_port);
   U201 : NAND2_X1 port map( A1 => n119, A2 => n171_port, ZN => n125);
   U202 : NAND2_X1 port map( A1 => n153_port, A2 => n145_port, ZN => n136);
   U203 : INV_X1 port map( A => n119, ZN => n174_port);
   U204 : NAND2_X1 port map( A1 => n146_port, A2 => n145_port, ZN => n144_port)
                           ;
   U205 : INV_X1 port map( A => n145_port, ZN => n161_port);
   U206 : NAND2_X1 port map( A1 => n129, A2 => n130, ZN => n48);
   U207 : NAND2_X1 port map( A1 => n167_port, A2 => n133, ZN => n123);
   U208 : INV_X1 port map( A => n150_port, ZN => n173_port);
   U209 : NAND2_X1 port map( A1 => n110, A2 => n111, ZN => N145);
   U210 : NAND2_X1 port map( A1 => OUTPUT1_3_port, A2 => n13, ZN => n110);
   U211 : AOI22_X1 port map( A1 => OUTPUT2_3_port, A2 => n10, B1 => 
                           OUTPUT4_3_port, B2 => n7, ZN => n111);
   U212 : NAND2_X1 port map( A1 => n112, A2 => n113, ZN => N144);
   U213 : NAND2_X1 port map( A1 => OUTPUT1_2_port, A2 => n13, ZN => n112);
   U214 : AOI22_X1 port map( A1 => OUTPUT2_2_port, A2 => n10, B1 => 
                           OUTPUT4_2_port, B2 => n7, ZN => n113);
   U215 : NAND2_X1 port map( A1 => n114, A2 => n115, ZN => N143);
   U216 : NAND2_X1 port map( A1 => OUTPUT1_1_port, A2 => n13, ZN => n114);
   U217 : AOI22_X1 port map( A1 => OUTPUT2_1_port, A2 => n10, B1 => 
                           OUTPUT4_1_port, B2 => n7, ZN => n115);
   U218 : NOR2_X1 port map( A1 => FUNC(0), A2 => FUNC(1), ZN => n147_port);
   U219 : OAI211_X1 port map( C1 => n126, C2 => n127, A => n128, B => n48, ZN 
                           => N206);
   U220 : OAI21_X1 port map( B1 => n131, B2 => n130, A => n174_port, ZN => n128
                           );
   U224 : NOR3_X1 port map( A1 => n169_port, A2 => FUNC(2), A3 => n161_port, ZN
                           => n131);
   U225 : NOR2_X1 port map( A1 => n166_port, A2 => FUNC(1), ZN => n145_port);
   U226 : NOR2_X1 port map( A1 => n168_port, A2 => FUNC(3), ZN => n146_port);
   U227 : NAND2_X1 port map( A1 => FUNC(5), A2 => n172_port, ZN => n127);
   U228 : NAND2_X1 port map( A1 => FUNC(5), A2 => FUNC(4), ZN => n119);
   U229 : INV_X1 port map( A => FUNC(3), ZN => n169_port);
   U230 : INV_X1 port map( A => FUNC(2), ZN => n168_port);
   U231 : NOR2_X1 port map( A1 => FUNC(4), A2 => FUNC(5), ZN => n150_port);
   U232 : NOR2_X1 port map( A1 => n172_port, A2 => FUNC(5), ZN => n129);
   U233 : INV_X1 port map( A => FUNC(0), ZN => n166_port);
   U234 : INV_X1 port map( A => FUNC(4), ZN => n172_port);
   U235 : AND2_X1 port map( A1 => FUNC(1), A2 => n166_port, ZN => n133);
   U236 : INV_X1 port map( A => DATA2(3), ZN => n27);
   U237 : NAND2_X1 port map( A1 => n116, A2 => n117, ZN => N142);
   U238 : AOI22_X1 port map( A1 => OUTPUT3_0_port, A2 => n55, B1 => 
                           OUTPUT1_0_port, B2 => n15, ZN => n116);
   U239 : AOI22_X1 port map( A1 => OUTPUT2_0_port, A2 => n10, B1 => 
                           OUTPUT4_0_port, B2 => n7, ZN => n117);
   U240 : INV_X1 port map( A => DATA2(0), ZN => n22);
   U241 : INV_X1 port map( A => DATA2(1), ZN => n23);
   U242 : INV_X1 port map( A => n25, ZN => n24);
   U243 : INV_X1 port map( A => DATA2(2), ZN => n25);
   U244 : INV_X1 port map( A => DATA2(4), ZN => n28);

end SYN_Architectural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity regFFD_NBIT6_0 is

   port( CK, RESET, ENABLE : in std_logic;  D : in std_logic_vector (5 downto 
         0);  Q : out std_logic_vector (5 downto 0));

end regFFD_NBIT6_0;

architecture SYN_ASYNCHBEHAV of regFFD_NBIT6_0 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      , n17, n18 : std_logic;

begin
   
   Q_reg_5_inst : DFFR_X1 port map( D => n18, CK => CK, RN => RESET, Q => Q(5),
                           QN => n12);
   Q_reg_2_inst : DFFR_X1 port map( D => n15, CK => CK, RN => RESET, Q => Q(2),
                           QN => n9);
   Q_reg_1_inst : DFFR_X1 port map( D => n14, CK => CK, RN => RESET, Q => Q(1),
                           QN => n8);
   Q_reg_0_inst : DFFR_X1 port map( D => n13, CK => CK, RN => RESET, Q => Q(0),
                           QN => n7);
   Q_reg_3_inst : DFFR_X1 port map( D => n16, CK => CK, RN => RESET, Q => Q(3),
                           QN => n10);
   Q_reg_4_inst : DFFR_X1 port map( D => n17, CK => CK, RN => RESET, Q => Q(4),
                           QN => n11);
   U2 : OAI21_X1 port map( B1 => n9, B2 => ENABLE, A => n3, ZN => n15);
   U3 : NAND2_X1 port map( A1 => D(2), A2 => ENABLE, ZN => n3);
   U4 : OAI21_X1 port map( B1 => n8, B2 => ENABLE, A => n2, ZN => n14);
   U5 : NAND2_X1 port map( A1 => D(1), A2 => ENABLE, ZN => n2);
   U6 : OAI21_X1 port map( B1 => n7, B2 => ENABLE, A => n1, ZN => n13);
   U7 : NAND2_X1 port map( A1 => ENABLE, A2 => D(0), ZN => n1);
   U8 : OAI21_X1 port map( B1 => n12, B2 => ENABLE, A => n6, ZN => n18);
   U9 : NAND2_X1 port map( A1 => D(5), A2 => ENABLE, ZN => n6);
   U10 : OAI21_X1 port map( B1 => n11, B2 => ENABLE, A => n5, ZN => n17);
   U11 : NAND2_X1 port map( A1 => D(4), A2 => ENABLE, ZN => n5);
   U12 : OAI21_X1 port map( B1 => n10, B2 => ENABLE, A => n4, ZN => n16);
   U13 : NAND2_X1 port map( A1 => D(3), A2 => ENABLE, ZN => n4);

end SYN_ASYNCHBEHAV;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity regFFD_NBIT5_0 is

   port( CK, RESET, ENABLE : in std_logic;  D : in std_logic_vector (4 downto 
         0);  Q : out std_logic_vector (4 downto 0));

end regFFD_NBIT5_0;

architecture SYN_ASYNCHBEHAV of regFFD_NBIT5_0 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15 : 
      std_logic;

begin
   
   Q_reg_2_inst : DFFR_X1 port map( D => n13, CK => CK, RN => RESET, Q => Q(2),
                           QN => n8);
   Q_reg_3_inst : DFFR_X1 port map( D => n14, CK => CK, RN => RESET, Q => Q(3),
                           QN => n9);
   Q_reg_0_inst : DFFR_X1 port map( D => n11, CK => CK, RN => RESET, Q => Q(0),
                           QN => n6);
   Q_reg_4_inst : DFFR_X1 port map( D => n15, CK => CK, RN => RESET, Q => Q(4),
                           QN => n10);
   Q_reg_1_inst : DFFR_X1 port map( D => n12, CK => CK, RN => RESET, Q => Q(1),
                           QN => n7);
   U2 : OAI21_X1 port map( B1 => n7, B2 => ENABLE, A => n2, ZN => n12);
   U3 : NAND2_X1 port map( A1 => D(1), A2 => ENABLE, ZN => n2);
   U4 : OAI21_X1 port map( B1 => n8, B2 => ENABLE, A => n3, ZN => n13);
   U5 : NAND2_X1 port map( A1 => D(2), A2 => ENABLE, ZN => n3);
   U6 : OAI21_X1 port map( B1 => n9, B2 => ENABLE, A => n4, ZN => n14);
   U7 : NAND2_X1 port map( A1 => D(3), A2 => ENABLE, ZN => n4);
   U8 : OAI21_X1 port map( B1 => n10, B2 => ENABLE, A => n5, ZN => n15);
   U9 : NAND2_X1 port map( A1 => D(4), A2 => ENABLE, ZN => n5);
   U10 : OAI21_X1 port map( B1 => n6, B2 => ENABLE, A => n1, ZN => n11);
   U11 : NAND2_X1 port map( A1 => ENABLE, A2 => D(0), ZN => n1);

end SYN_ASYNCHBEHAV;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FF_0 is

   port( CLK, RESET, EN, D : in std_logic;  Q : out std_logic);

end FF_0;

architecture SYN_SYNC_BHV of FF_0 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n3, n4, n1, n2, n_1152 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFF_X1 port map( D => n4, CK => CLK, Q => Q_port, QN => n_1152);
   U3 : NOR2_X1 port map( A1 => n3, A2 => n1, ZN => n4);
   U4 : AOI22_X1 port map( A1 => EN, A2 => D, B1 => Q_port, B2 => n2, ZN => n3)
                           ;
   U5 : INV_X1 port map( A => EN, ZN => n2);
   U6 : INV_X1 port map( A => RESET, ZN => n1);

end SYN_SYNC_BHV;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity windRF_M8_N8_F5_NBIT32 is

   port( CLK, RESET, ENABLE, CALL, RETRN : in std_logic;  FILL, SPILL : out 
         std_logic;  BUSin : in std_logic_vector (31 downto 0);  BUSout : out 
         std_logic_vector (31 downto 0);  RD1, RD2, WR : in std_logic;  ADD_WR,
         ADD_RD1, ADD_RD2 : in std_logic_vector (4 downto 0);  DATAIN : in 
         std_logic_vector (31 downto 0);  OUT1, OUT2 : out std_logic_vector (31
         downto 0);  wr_signal : in std_logic);

end windRF_M8_N8_F5_NBIT32;

architecture SYN_bhv of windRF_M8_N8_F5_NBIT32 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component windRF_M8_N8_F5_NBIT32_DW01_add_5
      port( A, B : in std_logic_vector (6 downto 0);  CI : in std_logic;  SUM :
            out std_logic_vector (6 downto 0);  CO : out std_logic);
   end component;
   
   component windRF_M8_N8_F5_NBIT32_DW01_add_3
      port( A, B : in std_logic_vector (6 downto 0);  CI : in std_logic;  SUM :
            out std_logic_vector (6 downto 0);  CO : out std_logic);
   end component;
   
   component windRF_M8_N8_F5_NBIT32_DW01_add_1
      port( A, B : in std_logic_vector (6 downto 0);  CI : in std_logic;  SUM :
            out std_logic_vector (6 downto 0);  CO : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal REGISTERS_11_31_port, REGISTERS_11_30_port, REGISTERS_11_29_port, 
      REGISTERS_11_28_port, REGISTERS_11_27_port, REGISTERS_11_26_port, 
      REGISTERS_11_25_port, REGISTERS_11_24_port, REGISTERS_11_23_port, 
      REGISTERS_11_22_port, REGISTERS_11_21_port, REGISTERS_11_20_port, 
      REGISTERS_11_19_port, REGISTERS_11_18_port, REGISTERS_11_17_port, 
      REGISTERS_11_16_port, REGISTERS_11_15_port, REGISTERS_11_14_port, 
      REGISTERS_11_13_port, REGISTERS_11_12_port, REGISTERS_11_11_port, 
      REGISTERS_11_10_port, REGISTERS_11_9_port, REGISTERS_11_8_port, 
      REGISTERS_11_7_port, REGISTERS_11_6_port, REGISTERS_11_5_port, 
      REGISTERS_11_4_port, REGISTERS_11_3_port, REGISTERS_11_2_port, 
      REGISTERS_11_1_port, REGISTERS_11_0_port, REGISTERS_12_31_port, 
      REGISTERS_12_30_port, REGISTERS_12_29_port, REGISTERS_12_28_port, 
      REGISTERS_12_27_port, REGISTERS_12_26_port, REGISTERS_12_25_port, 
      REGISTERS_12_24_port, REGISTERS_12_23_port, REGISTERS_12_22_port, 
      REGISTERS_12_21_port, REGISTERS_12_20_port, REGISTERS_12_19_port, 
      REGISTERS_12_18_port, REGISTERS_12_17_port, REGISTERS_12_16_port, 
      REGISTERS_12_15_port, REGISTERS_12_14_port, REGISTERS_12_13_port, 
      REGISTERS_12_12_port, REGISTERS_12_11_port, REGISTERS_12_10_port, 
      REGISTERS_12_9_port, REGISTERS_12_8_port, REGISTERS_12_7_port, 
      REGISTERS_12_6_port, REGISTERS_12_5_port, REGISTERS_12_4_port, 
      REGISTERS_12_3_port, REGISTERS_12_2_port, REGISTERS_12_1_port, 
      REGISTERS_12_0_port, REGISTERS_16_31_port, REGISTERS_16_30_port, 
      REGISTERS_16_29_port, REGISTERS_16_28_port, REGISTERS_16_27_port, 
      REGISTERS_16_26_port, REGISTERS_16_25_port, REGISTERS_16_24_port, 
      REGISTERS_16_23_port, REGISTERS_16_22_port, REGISTERS_16_21_port, 
      REGISTERS_16_20_port, REGISTERS_16_19_port, REGISTERS_16_18_port, 
      REGISTERS_16_17_port, REGISTERS_16_16_port, REGISTERS_16_15_port, 
      REGISTERS_16_14_port, REGISTERS_16_13_port, REGISTERS_16_12_port, 
      REGISTERS_16_11_port, REGISTERS_16_10_port, REGISTERS_16_9_port, 
      REGISTERS_16_8_port, REGISTERS_16_7_port, REGISTERS_16_6_port, 
      REGISTERS_16_5_port, REGISTERS_16_4_port, REGISTERS_16_3_port, 
      REGISTERS_16_2_port, REGISTERS_16_1_port, REGISTERS_16_0_port, 
      REGISTERS_17_31_port, REGISTERS_17_30_port, REGISTERS_17_29_port, 
      REGISTERS_17_28_port, REGISTERS_17_27_port, REGISTERS_17_26_port, 
      REGISTERS_17_25_port, REGISTERS_17_24_port, REGISTERS_17_23_port, 
      REGISTERS_17_22_port, REGISTERS_17_21_port, REGISTERS_17_20_port, 
      REGISTERS_17_19_port, REGISTERS_17_18_port, REGISTERS_17_17_port, 
      REGISTERS_17_16_port, REGISTERS_17_15_port, REGISTERS_17_14_port, 
      REGISTERS_17_13_port, REGISTERS_17_12_port, REGISTERS_17_11_port, 
      REGISTERS_17_10_port, REGISTERS_17_9_port, REGISTERS_17_8_port, 
      REGISTERS_17_7_port, REGISTERS_17_6_port, REGISTERS_17_5_port, 
      REGISTERS_17_4_port, REGISTERS_17_3_port, REGISTERS_17_2_port, 
      REGISTERS_17_1_port, REGISTERS_17_0_port, REGISTERS_18_31_port, 
      REGISTERS_18_30_port, REGISTERS_18_29_port, REGISTERS_18_28_port, 
      REGISTERS_18_27_port, REGISTERS_18_26_port, REGISTERS_18_25_port, 
      REGISTERS_18_24_port, REGISTERS_18_23_port, REGISTERS_18_22_port, 
      REGISTERS_18_21_port, REGISTERS_18_20_port, REGISTERS_18_19_port, 
      REGISTERS_18_18_port, REGISTERS_18_17_port, REGISTERS_18_16_port, 
      REGISTERS_18_15_port, REGISTERS_18_14_port, REGISTERS_18_13_port, 
      REGISTERS_18_12_port, REGISTERS_18_11_port, REGISTERS_18_10_port, 
      REGISTERS_18_9_port, REGISTERS_18_8_port, REGISTERS_18_7_port, 
      REGISTERS_18_6_port, REGISTERS_18_5_port, REGISTERS_18_4_port, 
      REGISTERS_18_3_port, REGISTERS_18_2_port, REGISTERS_18_1_port, 
      REGISTERS_18_0_port, REGISTERS_19_31_port, REGISTERS_19_30_port, 
      REGISTERS_19_29_port, REGISTERS_19_28_port, REGISTERS_19_27_port, 
      REGISTERS_19_26_port, REGISTERS_19_25_port, REGISTERS_19_24_port, 
      REGISTERS_19_23_port, REGISTERS_19_22_port, REGISTERS_19_21_port, 
      REGISTERS_19_20_port, REGISTERS_19_19_port, REGISTERS_19_18_port, 
      REGISTERS_19_17_port, REGISTERS_19_16_port, REGISTERS_19_15_port, 
      REGISTERS_19_14_port, REGISTERS_19_13_port, REGISTERS_19_12_port, 
      REGISTERS_19_11_port, REGISTERS_19_10_port, REGISTERS_19_9_port, 
      REGISTERS_19_8_port, REGISTERS_19_7_port, REGISTERS_19_6_port, 
      REGISTERS_19_5_port, REGISTERS_19_4_port, REGISTERS_19_3_port, 
      REGISTERS_19_2_port, REGISTERS_19_1_port, REGISTERS_19_0_port, 
      REGISTERS_20_31_port, REGISTERS_20_30_port, REGISTERS_20_29_port, 
      REGISTERS_20_28_port, REGISTERS_20_27_port, REGISTERS_20_26_port, 
      REGISTERS_20_25_port, REGISTERS_20_24_port, REGISTERS_20_23_port, 
      REGISTERS_20_22_port, REGISTERS_20_21_port, REGISTERS_20_20_port, 
      REGISTERS_20_19_port, REGISTERS_20_18_port, REGISTERS_20_17_port, 
      REGISTERS_20_16_port, REGISTERS_20_15_port, REGISTERS_20_14_port, 
      REGISTERS_20_13_port, REGISTERS_20_12_port, REGISTERS_20_11_port, 
      REGISTERS_20_10_port, REGISTERS_20_9_port, REGISTERS_20_8_port, 
      REGISTERS_20_7_port, REGISTERS_20_6_port, REGISTERS_20_5_port, 
      REGISTERS_20_4_port, REGISTERS_20_3_port, REGISTERS_20_2_port, 
      REGISTERS_20_1_port, REGISTERS_20_0_port, REGISTERS_21_31_port, 
      REGISTERS_21_30_port, REGISTERS_21_29_port, REGISTERS_21_28_port, 
      REGISTERS_21_27_port, REGISTERS_21_26_port, REGISTERS_21_25_port, 
      REGISTERS_21_24_port, REGISTERS_21_23_port, REGISTERS_21_22_port, 
      REGISTERS_21_21_port, REGISTERS_21_20_port, REGISTERS_21_19_port, 
      REGISTERS_21_18_port, REGISTERS_21_17_port, REGISTERS_21_16_port, 
      REGISTERS_21_15_port, REGISTERS_21_14_port, REGISTERS_21_13_port, 
      REGISTERS_21_12_port, REGISTERS_21_11_port, REGISTERS_21_10_port, 
      REGISTERS_21_9_port, REGISTERS_21_8_port, REGISTERS_21_7_port, 
      REGISTERS_21_6_port, REGISTERS_21_5_port, REGISTERS_21_4_port, 
      REGISTERS_21_3_port, REGISTERS_21_2_port, REGISTERS_21_1_port, 
      REGISTERS_21_0_port, REGISTERS_33_31_port, REGISTERS_33_30_port, 
      REGISTERS_33_29_port, REGISTERS_33_28_port, REGISTERS_33_27_port, 
      REGISTERS_33_26_port, REGISTERS_33_25_port, REGISTERS_33_24_port, 
      REGISTERS_33_23_port, REGISTERS_33_22_port, REGISTERS_33_21_port, 
      REGISTERS_33_20_port, REGISTERS_33_19_port, REGISTERS_33_18_port, 
      REGISTERS_33_17_port, REGISTERS_33_16_port, REGISTERS_33_15_port, 
      REGISTERS_33_14_port, REGISTERS_33_13_port, REGISTERS_33_12_port, 
      REGISTERS_33_11_port, REGISTERS_33_10_port, REGISTERS_33_9_port, 
      REGISTERS_33_8_port, REGISTERS_33_7_port, REGISTERS_33_6_port, 
      REGISTERS_33_5_port, REGISTERS_33_4_port, REGISTERS_33_3_port, 
      REGISTERS_33_2_port, REGISTERS_33_1_port, REGISTERS_33_0_port, 
      REGISTERS_34_31_port, REGISTERS_34_30_port, REGISTERS_34_29_port, 
      REGISTERS_34_28_port, REGISTERS_34_27_port, REGISTERS_34_26_port, 
      REGISTERS_34_25_port, REGISTERS_34_24_port, REGISTERS_34_23_port, 
      REGISTERS_34_22_port, REGISTERS_34_21_port, REGISTERS_34_20_port, 
      REGISTERS_34_19_port, REGISTERS_34_18_port, REGISTERS_34_17_port, 
      REGISTERS_34_16_port, REGISTERS_34_15_port, REGISTERS_34_14_port, 
      REGISTERS_34_13_port, REGISTERS_34_12_port, REGISTERS_34_11_port, 
      REGISTERS_34_10_port, REGISTERS_34_9_port, REGISTERS_34_8_port, 
      REGISTERS_34_7_port, REGISTERS_34_6_port, REGISTERS_34_5_port, 
      REGISTERS_34_4_port, REGISTERS_34_3_port, REGISTERS_34_2_port, 
      REGISTERS_34_1_port, REGISTERS_34_0_port, REGISTERS_38_31_port, 
      REGISTERS_38_30_port, REGISTERS_38_29_port, REGISTERS_38_28_port, 
      REGISTERS_38_27_port, REGISTERS_38_26_port, REGISTERS_38_25_port, 
      REGISTERS_38_24_port, REGISTERS_38_23_port, REGISTERS_38_22_port, 
      REGISTERS_38_21_port, REGISTERS_38_20_port, REGISTERS_38_19_port, 
      REGISTERS_38_18_port, REGISTERS_38_17_port, REGISTERS_38_16_port, 
      REGISTERS_38_15_port, REGISTERS_38_14_port, REGISTERS_38_13_port, 
      REGISTERS_38_12_port, REGISTERS_38_11_port, REGISTERS_38_10_port, 
      REGISTERS_38_9_port, REGISTERS_38_8_port, REGISTERS_38_7_port, 
      REGISTERS_38_6_port, REGISTERS_38_5_port, REGISTERS_38_4_port, 
      REGISTERS_38_3_port, REGISTERS_38_2_port, REGISTERS_38_1_port, 
      REGISTERS_38_0_port, REGISTERS_39_31_port, REGISTERS_39_30_port, 
      REGISTERS_39_29_port, REGISTERS_39_28_port, REGISTERS_39_27_port, 
      REGISTERS_39_26_port, REGISTERS_39_25_port, REGISTERS_39_24_port, 
      REGISTERS_39_23_port, REGISTERS_39_22_port, REGISTERS_39_21_port, 
      REGISTERS_39_20_port, REGISTERS_39_19_port, REGISTERS_39_18_port, 
      REGISTERS_39_17_port, REGISTERS_39_16_port, REGISTERS_39_15_port, 
      REGISTERS_39_14_port, REGISTERS_39_13_port, REGISTERS_39_12_port, 
      REGISTERS_39_11_port, REGISTERS_39_10_port, REGISTERS_39_9_port, 
      REGISTERS_39_8_port, REGISTERS_39_7_port, REGISTERS_39_6_port, 
      REGISTERS_39_5_port, REGISTERS_39_4_port, REGISTERS_39_3_port, 
      REGISTERS_39_2_port, REGISTERS_39_1_port, REGISTERS_39_0_port, 
      REGISTERS_40_31_port, REGISTERS_40_30_port, REGISTERS_40_29_port, 
      REGISTERS_40_28_port, REGISTERS_40_27_port, REGISTERS_40_26_port, 
      REGISTERS_40_25_port, REGISTERS_40_24_port, REGISTERS_40_23_port, 
      REGISTERS_40_22_port, REGISTERS_40_21_port, REGISTERS_40_20_port, 
      REGISTERS_40_19_port, REGISTERS_40_18_port, REGISTERS_40_17_port, 
      REGISTERS_40_16_port, REGISTERS_40_15_port, REGISTERS_40_14_port, 
      REGISTERS_40_13_port, REGISTERS_40_12_port, REGISTERS_40_11_port, 
      REGISTERS_40_10_port, REGISTERS_40_9_port, REGISTERS_40_8_port, 
      REGISTERS_40_7_port, REGISTERS_40_6_port, REGISTERS_40_5_port, 
      REGISTERS_40_4_port, REGISTERS_40_3_port, REGISTERS_40_2_port, 
      REGISTERS_40_1_port, REGISTERS_40_0_port, REGISTERS_41_31_port, 
      REGISTERS_41_30_port, REGISTERS_41_29_port, REGISTERS_41_28_port, 
      REGISTERS_41_27_port, REGISTERS_41_26_port, REGISTERS_41_25_port, 
      REGISTERS_41_24_port, REGISTERS_41_23_port, REGISTERS_41_22_port, 
      REGISTERS_41_21_port, REGISTERS_41_20_port, REGISTERS_41_19_port, 
      REGISTERS_41_18_port, REGISTERS_41_17_port, REGISTERS_41_16_port, 
      REGISTERS_41_15_port, REGISTERS_41_14_port, REGISTERS_41_13_port, 
      REGISTERS_41_12_port, REGISTERS_41_11_port, REGISTERS_41_10_port, 
      REGISTERS_41_9_port, REGISTERS_41_8_port, REGISTERS_41_7_port, 
      REGISTERS_41_6_port, REGISTERS_41_5_port, REGISTERS_41_4_port, 
      REGISTERS_41_3_port, REGISTERS_41_2_port, REGISTERS_41_1_port, 
      REGISTERS_41_0_port, REGISTERS_42_31_port, REGISTERS_42_30_port, 
      REGISTERS_42_29_port, REGISTERS_42_28_port, REGISTERS_42_27_port, 
      REGISTERS_42_26_port, REGISTERS_42_25_port, REGISTERS_42_24_port, 
      REGISTERS_42_23_port, REGISTERS_42_22_port, REGISTERS_42_21_port, 
      REGISTERS_42_20_port, REGISTERS_42_19_port, REGISTERS_42_18_port, 
      REGISTERS_42_17_port, REGISTERS_42_16_port, REGISTERS_42_15_port, 
      REGISTERS_42_14_port, REGISTERS_42_13_port, REGISTERS_42_12_port, 
      REGISTERS_42_11_port, REGISTERS_42_10_port, REGISTERS_42_9_port, 
      REGISTERS_42_8_port, REGISTERS_42_7_port, REGISTERS_42_6_port, 
      REGISTERS_42_5_port, REGISTERS_42_4_port, REGISTERS_42_3_port, 
      REGISTERS_42_2_port, REGISTERS_42_1_port, REGISTERS_42_0_port, 
      REGISTERS_43_31_port, REGISTERS_43_30_port, REGISTERS_43_29_port, 
      REGISTERS_43_28_port, REGISTERS_43_27_port, REGISTERS_43_26_port, 
      REGISTERS_43_25_port, REGISTERS_43_24_port, REGISTERS_43_23_port, 
      REGISTERS_43_22_port, REGISTERS_43_21_port, REGISTERS_43_20_port, 
      REGISTERS_43_19_port, REGISTERS_43_18_port, REGISTERS_43_17_port, 
      REGISTERS_43_16_port, REGISTERS_43_15_port, REGISTERS_43_14_port, 
      REGISTERS_43_13_port, REGISTERS_43_12_port, REGISTERS_43_11_port, 
      REGISTERS_43_10_port, REGISTERS_43_9_port, REGISTERS_43_8_port, 
      REGISTERS_43_7_port, REGISTERS_43_6_port, REGISTERS_43_5_port, 
      REGISTERS_43_4_port, REGISTERS_43_3_port, REGISTERS_43_2_port, 
      REGISTERS_43_1_port, REGISTERS_43_0_port, REGISTERS_44_31_port, 
      REGISTERS_44_30_port, REGISTERS_44_29_port, REGISTERS_44_28_port, 
      REGISTERS_44_27_port, REGISTERS_44_26_port, REGISTERS_44_25_port, 
      REGISTERS_44_24_port, REGISTERS_44_23_port, REGISTERS_44_22_port, 
      REGISTERS_44_21_port, REGISTERS_44_20_port, REGISTERS_44_19_port, 
      REGISTERS_44_18_port, REGISTERS_44_17_port, REGISTERS_44_16_port, 
      REGISTERS_44_15_port, REGISTERS_44_14_port, REGISTERS_44_13_port, 
      REGISTERS_44_12_port, REGISTERS_44_11_port, REGISTERS_44_10_port, 
      REGISTERS_44_9_port, REGISTERS_44_8_port, REGISTERS_44_7_port, 
      REGISTERS_44_6_port, REGISTERS_44_5_port, REGISTERS_44_4_port, 
      REGISTERS_44_3_port, REGISTERS_44_2_port, REGISTERS_44_1_port, 
      REGISTERS_44_0_port, REGISTERS_45_31_port, REGISTERS_45_30_port, 
      REGISTERS_45_29_port, REGISTERS_45_28_port, REGISTERS_45_27_port, 
      REGISTERS_45_26_port, REGISTERS_45_25_port, REGISTERS_45_24_port, 
      REGISTERS_45_23_port, REGISTERS_45_22_port, REGISTERS_45_21_port, 
      REGISTERS_45_20_port, REGISTERS_45_19_port, REGISTERS_45_18_port, 
      REGISTERS_45_17_port, REGISTERS_45_16_port, REGISTERS_45_15_port, 
      REGISTERS_45_14_port, REGISTERS_45_13_port, REGISTERS_45_12_port, 
      REGISTERS_45_11_port, REGISTERS_45_10_port, REGISTERS_45_9_port, 
      REGISTERS_45_8_port, REGISTERS_45_7_port, REGISTERS_45_6_port, 
      REGISTERS_45_5_port, REGISTERS_45_4_port, REGISTERS_45_3_port, 
      REGISTERS_45_2_port, REGISTERS_45_1_port, REGISTERS_45_0_port, 
      REGISTERS_49_31_port, REGISTERS_49_30_port, REGISTERS_49_29_port, 
      REGISTERS_49_28_port, REGISTERS_49_27_port, REGISTERS_49_26_port, 
      REGISTERS_49_25_port, REGISTERS_49_24_port, REGISTERS_49_23_port, 
      REGISTERS_49_22_port, REGISTERS_49_21_port, REGISTERS_49_20_port, 
      REGISTERS_49_19_port, REGISTERS_49_18_port, REGISTERS_49_17_port, 
      REGISTERS_49_16_port, REGISTERS_49_15_port, REGISTERS_49_14_port, 
      REGISTERS_49_13_port, REGISTERS_49_12_port, REGISTERS_49_11_port, 
      REGISTERS_49_10_port, REGISTERS_49_9_port, REGISTERS_49_8_port, 
      REGISTERS_49_7_port, REGISTERS_49_6_port, REGISTERS_49_5_port, 
      REGISTERS_49_4_port, REGISTERS_49_3_port, REGISTERS_49_2_port, 
      REGISTERS_49_1_port, REGISTERS_49_0_port, REGISTERS_50_31_port, 
      REGISTERS_50_30_port, REGISTERS_50_29_port, REGISTERS_50_28_port, 
      REGISTERS_50_27_port, REGISTERS_50_26_port, REGISTERS_50_25_port, 
      REGISTERS_50_24_port, REGISTERS_50_23_port, REGISTERS_50_22_port, 
      REGISTERS_50_21_port, REGISTERS_50_20_port, REGISTERS_50_19_port, 
      REGISTERS_50_18_port, REGISTERS_50_17_port, REGISTERS_50_16_port, 
      REGISTERS_50_15_port, REGISTERS_50_14_port, REGISTERS_50_13_port, 
      REGISTERS_50_12_port, REGISTERS_50_11_port, REGISTERS_50_10_port, 
      REGISTERS_50_9_port, REGISTERS_50_8_port, REGISTERS_50_7_port, 
      REGISTERS_50_6_port, REGISTERS_50_5_port, REGISTERS_50_4_port, 
      REGISTERS_50_3_port, REGISTERS_50_2_port, REGISTERS_50_1_port, 
      REGISTERS_50_0_port, REGISTERS_51_31_port, REGISTERS_51_30_port, 
      REGISTERS_51_29_port, REGISTERS_51_28_port, REGISTERS_51_27_port, 
      REGISTERS_51_26_port, REGISTERS_51_25_port, REGISTERS_51_24_port, 
      REGISTERS_51_23_port, REGISTERS_51_22_port, REGISTERS_51_21_port, 
      REGISTERS_51_20_port, REGISTERS_51_19_port, REGISTERS_51_18_port, 
      REGISTERS_51_17_port, REGISTERS_51_16_port, REGISTERS_51_15_port, 
      REGISTERS_51_14_port, REGISTERS_51_13_port, REGISTERS_51_12_port, 
      REGISTERS_51_11_port, REGISTERS_51_10_port, REGISTERS_51_9_port, 
      REGISTERS_51_8_port, REGISTERS_51_7_port, REGISTERS_51_6_port, 
      REGISTERS_51_5_port, REGISTERS_51_4_port, REGISTERS_51_3_port, 
      REGISTERS_51_2_port, REGISTERS_51_1_port, REGISTERS_51_0_port, 
      REGISTERS_52_31_port, REGISTERS_52_30_port, REGISTERS_52_29_port, 
      REGISTERS_52_28_port, REGISTERS_52_27_port, REGISTERS_52_26_port, 
      REGISTERS_52_25_port, REGISTERS_52_24_port, REGISTERS_52_23_port, 
      REGISTERS_52_22_port, REGISTERS_52_21_port, REGISTERS_52_20_port, 
      REGISTERS_52_19_port, REGISTERS_52_18_port, REGISTERS_52_17_port, 
      REGISTERS_52_16_port, REGISTERS_52_15_port, REGISTERS_52_14_port, 
      REGISTERS_52_13_port, REGISTERS_52_12_port, REGISTERS_52_11_port, 
      REGISTERS_52_10_port, REGISTERS_52_9_port, REGISTERS_52_8_port, 
      REGISTERS_52_7_port, REGISTERS_52_6_port, REGISTERS_52_5_port, 
      REGISTERS_52_4_port, REGISTERS_52_3_port, REGISTERS_52_2_port, 
      REGISTERS_52_1_port, REGISTERS_52_0_port, REGISTERS_53_31_port, 
      REGISTERS_53_30_port, REGISTERS_53_29_port, REGISTERS_53_28_port, 
      REGISTERS_53_27_port, REGISTERS_53_26_port, REGISTERS_53_25_port, 
      REGISTERS_53_24_port, REGISTERS_53_23_port, REGISTERS_53_22_port, 
      REGISTERS_53_21_port, REGISTERS_53_20_port, REGISTERS_53_19_port, 
      REGISTERS_53_18_port, REGISTERS_53_17_port, REGISTERS_53_16_port, 
      REGISTERS_53_15_port, REGISTERS_53_14_port, REGISTERS_53_13_port, 
      REGISTERS_53_12_port, REGISTERS_53_11_port, REGISTERS_53_10_port, 
      REGISTERS_53_9_port, REGISTERS_53_8_port, REGISTERS_53_7_port, 
      REGISTERS_53_6_port, REGISTERS_53_5_port, REGISTERS_53_4_port, 
      REGISTERS_53_3_port, REGISTERS_53_2_port, REGISTERS_53_1_port, 
      REGISTERS_53_0_port, REGISTERS_54_31_port, REGISTERS_54_30_port, 
      REGISTERS_54_29_port, REGISTERS_54_28_port, REGISTERS_54_27_port, 
      REGISTERS_54_26_port, REGISTERS_54_25_port, REGISTERS_54_24_port, 
      REGISTERS_54_23_port, REGISTERS_54_22_port, REGISTERS_54_21_port, 
      REGISTERS_54_20_port, REGISTERS_54_19_port, REGISTERS_54_18_port, 
      REGISTERS_54_17_port, REGISTERS_54_16_port, REGISTERS_54_15_port, 
      REGISTERS_54_14_port, REGISTERS_54_13_port, REGISTERS_54_12_port, 
      REGISTERS_54_11_port, REGISTERS_54_10_port, REGISTERS_54_9_port, 
      REGISTERS_54_8_port, REGISTERS_54_7_port, REGISTERS_54_6_port, 
      REGISTERS_54_5_port, REGISTERS_54_4_port, REGISTERS_54_3_port, 
      REGISTERS_54_2_port, REGISTERS_54_1_port, REGISTERS_54_0_port, 
      REGISTERS_77_31_port, REGISTERS_77_30_port, REGISTERS_77_29_port, 
      REGISTERS_77_28_port, REGISTERS_77_27_port, REGISTERS_77_26_port, 
      REGISTERS_77_25_port, REGISTERS_77_24_port, REGISTERS_77_23_port, 
      REGISTERS_77_22_port, REGISTERS_77_21_port, REGISTERS_77_20_port, 
      REGISTERS_77_19_port, REGISTERS_77_18_port, REGISTERS_77_17_port, 
      REGISTERS_77_16_port, REGISTERS_77_15_port, REGISTERS_77_14_port, 
      REGISTERS_77_13_port, REGISTERS_77_12_port, REGISTERS_77_11_port, 
      REGISTERS_77_10_port, REGISTERS_77_9_port, REGISTERS_77_8_port, 
      REGISTERS_77_7_port, REGISTERS_77_6_port, REGISTERS_77_5_port, 
      REGISTERS_77_4_port, REGISTERS_77_3_port, REGISTERS_77_2_port, 
      REGISTERS_77_1_port, REGISTERS_77_0_port, REGISTERS_78_31_port, 
      REGISTERS_78_30_port, REGISTERS_78_29_port, REGISTERS_78_28_port, 
      REGISTERS_78_27_port, REGISTERS_78_26_port, REGISTERS_78_25_port, 
      REGISTERS_78_24_port, REGISTERS_78_23_port, REGISTERS_78_22_port, 
      REGISTERS_78_21_port, REGISTERS_78_20_port, REGISTERS_78_19_port, 
      REGISTERS_78_18_port, REGISTERS_78_17_port, REGISTERS_78_16_port, 
      REGISTERS_78_15_port, REGISTERS_78_14_port, REGISTERS_78_13_port, 
      REGISTERS_78_12_port, REGISTERS_78_11_port, REGISTERS_78_10_port, 
      REGISTERS_78_9_port, REGISTERS_78_8_port, REGISTERS_78_7_port, 
      REGISTERS_78_6_port, REGISTERS_78_5_port, REGISTERS_78_4_port, 
      REGISTERS_78_3_port, REGISTERS_78_2_port, REGISTERS_78_1_port, 
      REGISTERS_78_0_port, REGISTERS_82_31_port, REGISTERS_82_30_port, 
      REGISTERS_82_29_port, REGISTERS_82_28_port, REGISTERS_82_27_port, 
      REGISTERS_82_26_port, REGISTERS_82_25_port, REGISTERS_82_24_port, 
      REGISTERS_82_23_port, REGISTERS_82_22_port, REGISTERS_82_21_port, 
      REGISTERS_82_20_port, REGISTERS_82_19_port, REGISTERS_82_18_port, 
      REGISTERS_82_17_port, REGISTERS_82_16_port, REGISTERS_82_15_port, 
      REGISTERS_82_14_port, REGISTERS_82_13_port, REGISTERS_82_12_port, 
      REGISTERS_82_11_port, REGISTERS_82_10_port, REGISTERS_82_9_port, 
      REGISTERS_82_8_port, REGISTERS_82_7_port, REGISTERS_82_6_port, 
      REGISTERS_82_5_port, REGISTERS_82_4_port, REGISTERS_82_3_port, 
      REGISTERS_82_2_port, REGISTERS_82_1_port, REGISTERS_82_0_port, 
      REGISTERS_83_31_port, REGISTERS_83_30_port, REGISTERS_83_29_port, 
      REGISTERS_83_28_port, REGISTERS_83_27_port, REGISTERS_83_26_port, 
      REGISTERS_83_25_port, REGISTERS_83_24_port, REGISTERS_83_23_port, 
      REGISTERS_83_22_port, REGISTERS_83_21_port, REGISTERS_83_20_port, 
      REGISTERS_83_19_port, REGISTERS_83_18_port, REGISTERS_83_17_port, 
      REGISTERS_83_16_port, REGISTERS_83_15_port, REGISTERS_83_14_port, 
      REGISTERS_83_13_port, REGISTERS_83_12_port, REGISTERS_83_11_port, 
      REGISTERS_83_10_port, REGISTERS_83_9_port, REGISTERS_83_8_port, 
      REGISTERS_83_7_port, REGISTERS_83_6_port, REGISTERS_83_5_port, 
      REGISTERS_83_4_port, REGISTERS_83_3_port, REGISTERS_83_2_port, 
      REGISTERS_83_1_port, REGISTERS_83_0_port, REGISTERS_84_31_port, 
      REGISTERS_84_30_port, REGISTERS_84_29_port, REGISTERS_84_28_port, 
      REGISTERS_84_27_port, REGISTERS_84_26_port, REGISTERS_84_25_port, 
      REGISTERS_84_24_port, REGISTERS_84_23_port, REGISTERS_84_22_port, 
      REGISTERS_84_21_port, REGISTERS_84_20_port, REGISTERS_84_19_port, 
      REGISTERS_84_18_port, REGISTERS_84_17_port, REGISTERS_84_16_port, 
      REGISTERS_84_15_port, REGISTERS_84_14_port, REGISTERS_84_13_port, 
      REGISTERS_84_12_port, REGISTERS_84_11_port, REGISTERS_84_10_port, 
      REGISTERS_84_9_port, REGISTERS_84_8_port, REGISTERS_84_7_port, 
      REGISTERS_84_6_port, REGISTERS_84_5_port, REGISTERS_84_4_port, 
      REGISTERS_84_3_port, REGISTERS_84_2_port, REGISTERS_84_1_port, 
      REGISTERS_84_0_port, REGISTERS_85_31_port, REGISTERS_85_30_port, 
      REGISTERS_85_29_port, REGISTERS_85_28_port, REGISTERS_85_27_port, 
      REGISTERS_85_26_port, REGISTERS_85_25_port, REGISTERS_85_24_port, 
      REGISTERS_85_23_port, REGISTERS_85_22_port, REGISTERS_85_21_port, 
      REGISTERS_85_20_port, REGISTERS_85_19_port, REGISTERS_85_18_port, 
      REGISTERS_85_17_port, REGISTERS_85_16_port, REGISTERS_85_15_port, 
      REGISTERS_85_14_port, REGISTERS_85_13_port, REGISTERS_85_12_port, 
      REGISTERS_85_11_port, REGISTERS_85_10_port, REGISTERS_85_9_port, 
      REGISTERS_85_8_port, REGISTERS_85_7_port, REGISTERS_85_6_port, 
      REGISTERS_85_5_port, REGISTERS_85_4_port, REGISTERS_85_3_port, 
      REGISTERS_85_2_port, REGISTERS_85_1_port, REGISTERS_85_0_port, 
      REGISTERS_86_31_port, REGISTERS_86_30_port, REGISTERS_86_29_port, 
      REGISTERS_86_28_port, REGISTERS_86_27_port, REGISTERS_86_26_port, 
      REGISTERS_86_25_port, REGISTERS_86_24_port, REGISTERS_86_23_port, 
      REGISTERS_86_22_port, REGISTERS_86_21_port, REGISTERS_86_20_port, 
      REGISTERS_86_19_port, REGISTERS_86_18_port, REGISTERS_86_17_port, 
      REGISTERS_86_16_port, REGISTERS_86_15_port, REGISTERS_86_14_port, 
      REGISTERS_86_13_port, REGISTERS_86_12_port, REGISTERS_86_11_port, 
      REGISTERS_86_10_port, REGISTERS_86_9_port, REGISTERS_86_8_port, 
      REGISTERS_86_7_port, REGISTERS_86_6_port, REGISTERS_86_5_port, 
      REGISTERS_86_4_port, REGISTERS_86_3_port, REGISTERS_86_2_port, 
      REGISTERS_86_1_port, REGISTERS_86_0_port, REGISTERS_87_31_port, 
      REGISTERS_87_30_port, REGISTERS_87_29_port, REGISTERS_87_28_port, 
      REGISTERS_87_27_port, REGISTERS_87_26_port, REGISTERS_87_25_port, 
      REGISTERS_87_24_port, REGISTERS_87_23_port, REGISTERS_87_22_port, 
      REGISTERS_87_21_port, REGISTERS_87_20_port, REGISTERS_87_19_port, 
      REGISTERS_87_18_port, REGISTERS_87_17_port, REGISTERS_87_16_port, 
      REGISTERS_87_15_port, REGISTERS_87_14_port, REGISTERS_87_13_port, 
      REGISTERS_87_12_port, REGISTERS_87_11_port, REGISTERS_87_10_port, 
      REGISTERS_87_9_port, REGISTERS_87_8_port, REGISTERS_87_7_port, 
      REGISTERS_87_6_port, REGISTERS_87_5_port, REGISTERS_87_4_port, 
      REGISTERS_87_3_port, REGISTERS_87_2_port, REGISTERS_87_1_port, 
      REGISTERS_87_0_port, CWP_6_port, CWP_5_port, CWP_4_port, N2151, N2153, 
      N2154, N2155, N2156, N2157, N2158, N2159, N2163, N2164, N2165, N2166, 
      N8415, N8417, N8418, N8419, N8420, N8421, N8422, N8423, N8427, N8428, 
      N8429, N8430, N8559, N8561, N8562, N8563, N8564, N8565, N8566, N8567, 
      N8571, N8572, N8573, N8574, N8702, N8703, N8704, N8705, N8706, N8707, 
      N8708, N8709, N8710, N8711, N8712, N8713, N8714, N8715, N8716, N8717, 
      N8718, N8719, N8720, N8721, N8722, N8723, N8724, N8725, N8726, N8727, 
      N8728, N8729, N8730, N8731, N8732, N8733, N8734, N8735, N8736, N8737, 
      N8738, N8739, N8740, N8741, N8742, N8743, N8744, N8745, N8746, N8747, 
      N8748, N8749, N8750, N8751, N8752, N8753, N8754, N8755, N8756, N8757, 
      N8758, N8759, N8760, N8761, N8762, N8763, N8764, N8765, N8766, N8767, 
      N8787, N8788, N8789, N8790, N8791, N8833, N8834, n7, n11, n17, n80, n81, 
      n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96
      , n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, 
      n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, 
      n121, n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, 
      n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, 
      n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, 
      n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, 
      n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, 
      n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, 
      n193, n194, n195, n196, n197, n198, n199, n200, n201, n202, n203, n204, 
      n205, n206, n207, n208, n209, n210, n211, n212, n213, n214, n215, n216, 
      n217, n218, n219, n220, n221, n222, n223, n224, n225, n226, n227, n228, 
      n229, n230, n231, n232, n233, n234, n235, n236, n237, n238, n239, n240, 
      n241, n242, n243, n244, n245, n246, n247, n248, n249, n250, n251, n252, 
      n253, n254, n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, 
      n265, n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276, 
      n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287, n288, 
      n289, n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, 
      n301, n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, 
      n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323, n324, 
      n325, n326, n327, n328, n329, n330, n331, n332, n333, n334, n335, n336, 
      n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, n347, n348, 
      n349, n350, n351, n352, n353, n354, n355, n356, n357, n358, n359, n360, 
      n361, n362, n363, n364, n365, n366, n367, n368, n369, n370, n371, n372, 
      n373, n374, n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, 
      n385, n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, 
      n397, n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, 
      n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, 
      n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n496, 
      n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, 
      n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, 
      n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, 
      n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, 
      n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, 
      n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, 
      n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, 
      n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, n784, 
      n785, n786, n787, n788, n789, n790, n791, n792, n793, n794, n795, n796, 
      n797, n798, n799, n800, n801, n802, n803, n804, n805, n806, n807, n808, 
      n809, n810, n811, n812, n813, n814, n815, n816, n817, n818, n819, n820, 
      n821, n822, n823, n824, n825, n826, n827, n828, n829, n830, n831, n832, 
      n833, n834, n835, n836, n837, n838, n839, n840, n841, n842, n843, n844, 
      n845, n846, n847, n848, n849, n850, n851, n852, n853, n854, n855, n856, 
      n857, n858, n859, n860, n861, n862, n863, n864, n865, n866, n867, n868, 
      n869, n870, n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, 
      n881, n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892, 
      n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903, n904, 
      n905, n906, n907, n908, n909, n910, n911, n912, n913, n914, n915, n916, 
      n917, n918, n919, n920, n921, n922, n923, n924, n925, n926, n927, n928, 
      n929, n930, n931, n932, n933, n934, n935, n936, n937, n938, n939, n940, 
      n941, n942, n943, n944, n945, n946, n947, n948, n949, n950, n951, n952, 
      n953, n954, n955, n956, n957, n958, n959, n960, n961, n962, n963, n964, 
      n965, n966, n967, n968, n969, n970, n971, n972, n973, n974, n975, n976, 
      n977, n978, n979, n980, n981, n982, n983, n984, n985, n986, n987, n988, 
      n989, n990, n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000, 
      n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, 
      n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, 
      n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, 
      n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, 
      n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, 
      n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, 
      n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, 
      n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, 
      n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, 
      n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, 
      n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, 
      n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, 
      n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, 
      n1131, n1132, n1133, n1134, n1135, n1200, n1201, n1202, n1203, n1204, 
      n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214, 
      n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224, 
      n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234, 
      n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244, 
      n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254, 
      n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264, 
      n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274, 
      n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284, 
      n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294, 
      n1295, n1552, n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560, 
      n1561, n1562, n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570, 
      n1571, n1572, n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580, 
      n1581, n1582, n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590, 
      n1591, n1592, n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600, 
      n1601, n1602, n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610, 
      n1611, n1612, n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620, 
      n1621, n1622, n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630, 
      n1631, n1632, n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640, 
      n1641, n1642, n1643, n1644, n1645, n1646, n1647, n1840, n1841, n1842, 
      n1843, n1844, n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852, 
      n1853, n1854, n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862, 
      n1863, n1864, n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872, 
      n1873, n1874, n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882, 
      n1883, n1884, n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892, 
      n1893, n1894, n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902, 
      n1903, n1904, n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912, 
      n1913, n1914, n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922, 
      n1923, n1924, n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932, 
      n1933, n1934, n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942, 
      n1943, n1944, n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952, 
      n1953, n1954, n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962, 
      n1963, n1964, n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972, 
      n1973, n1974, n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982, 
      n1983, n1984, n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992, 
      n1993, n1994, n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002, 
      n2003, n2004, n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012, 
      n2013, n2014, n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022, 
      n2023, n2024, n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032, 
      n2033, n2034, n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042, 
      n2043, n2044, n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052, 
      n2053, n2054, n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062, 
      n2063, n2064, n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072, 
      n2073, n2074, n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082, 
      n2083, n2084, n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092, 
      n2093, n2094, n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102, 
      n2103, n2104, n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112, 
      n2113, n2114, n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122, 
      n2123, n2124, n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132, 
      n2133, n2134, n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142, 
      n2143, n2144, n2145, n2146, n2147, n2148, n2149, n2150, n2151_port, n2152
      , n2153_port, n2154_port, n2155_port, n2156_port, n2157_port, n2158_port,
      n2159_port, n2160, n2161, n2162, n2163_port, n2164_port, n2165_port, 
      n2166_port, n2167, n2168, n2169, n2170, n2171, n2172, n2173, n2174, n2175
      , n2176, n2177, n2178, n2179, n2180, n2181, n2182, n2183, n2184, n2185, 
      n2186, n2187, n2188, n2189, n2190, n2191, n2192, n2193, n2194, n2195, 
      n2196, n2197, n2198, n2199, n2200, n2201, n2202, n2203, n2204, n2205, 
      n2206, n2207, n2208, n2209, n2210, n2211, n2212, n2213, n2214, n2215, 
      n2216, n2217, n2218, n2219, n2220, n2221, n2222, n2223, n2224, n2225, 
      n2226, n2227, n2228, n2229, n2230, n2231, n2232, n2233, n2234, n2235, 
      n2236, n2237, n2238, n2239, n2240, n2241, n2242, n2243, n2244, n2245, 
      n2246, n2247, n2248, n2249, n2250, n2251, n2252, n2253, n2254, n2255, 
      n2256, n2257, n2258, n2259, n2260, n2261, n2262, n2263, n2264, n2265, 
      n2266, n2267, n2268, n2269, n2270, n2271, n2272, n2273, n2274, n2275, 
      n2276, n2277, n2278, n2279, n2280, n2281, n2282, n2283, n2284, n2285, 
      n2286, n2287, n2288, n2289, n2290, n2291, n2292, n2293, n2294, n2295, 
      n2296, n2297, n2298, n2299, n2300, n2301, n2302, n2303, n2304, n2305, 
      n2306, n2307, n2308, n2309, n2310, n2311, n2312, n2313, n2314, n2315, 
      n2316, n2317, n2318, n2319, n2320, n2321, n2322, n2323, n2324, n2325, 
      n2326, n2327, n2328, n2329, n2330, n2331, n2332, n2333, n2334, n2335, 
      n2336, n2337, n2338, n2339, n2340, n2341, n2342, n2343, n2344, n2345, 
      n2346, n2347, n2348, n2349, n2350, n2351, n2352, n2353, n2354, n2355, 
      n2356, n2357, n2358, n2359, n2360, n2361, n2362, n2363, n2364, n2365, 
      n2366, n2367, n2368, n2369, n2370, n2371, n2372, n2373, n2374, n2375, 
      n2376, n2377, n2378, n2379, n2380, n2381, n2382, n2383, n2384, n2385, 
      n2386, n2387, n2388, n2389, n2390, n2391, n2392, n2393, n2394, n2395, 
      n2396, n2397, n2398, n2399, n2400, n2401, n2402, n2403, n2404, n2405, 
      n2406, n2407, n2408, n2409, n2410, n2411, n2412, n2413, n2414, n2415, 
      n2416, n2417, n2418, n2419, n2420, n2421, n2422, n2423, n2424, n2425, 
      n2426, n2427, n2428, n2429, n2430, n2431, n2432, n2433, n2434, n2435, 
      n2436, n2437, n2438, n2439, n2440, n2441, n2442, n2443, n2444, n2445, 
      n2446, n2447, n2448, n2449, n2450, n2451, n2452, n2453, n2454, n2455, 
      n2456, n2457, n2458, n2459, n2460, n2461, n2462, n2463, n2464, n2465, 
      n2466, n2467, n2468, n2469, n2470, n2471, n2472, n2473, n2474, n2475, 
      n2476, n2477, n2478, n2479, n2480, n2481, n2482, n2483, n2484, n2485, 
      n2486, n2487, n2488, n2489, n2490, n2491, n2492, n2493, n2494, n2495, 
      n2496, n2497, n2498, n2499, n2500, n2501, n2502, n2503, n2504, n2505, 
      n2506, n2507, n2508, n2509, n2510, n2511, n2512, n2513, n2514, n2515, 
      n2516, n2517, n2518, n2519, n2520, n2521, n2522, n2523, n2524, n2525, 
      n2526, n2527, n2528, n2529, n2530, n2531, n2532, n2533, n2534, n2535, 
      n2536, n2537, n2538, n2539, n2540, n2541, n2542, n2543, n2608, n2609, 
      n2610, n2611, n2612, n2613, n2614, n2615, n2616, n2617, n2618, n2619, 
      n2620, n2621, n2622, n2623, n2624, n2625, n2626, n2627, n2628, n2629, 
      n2630, n2631, n2632, n2633, n2634, n2635, n2636, n2637, n2638, n2639, 
      n2640, n2641, n2642, n2643, n2644, n2645, n2646, n2647, n2648, n2649, 
      n2650, n2651, n2652, n2653, n2654, n2655, n2656, n2657, n2658, n2659, 
      n2660, n2661, n2662, n2663, n2664, n2665, n2666, n2667, n2668, n2669, 
      n2670, n2671, n2672, n2673, n2674, n2675, n2676, n2677, n2678, n2679, 
      n2680, n2681, n2682, n2683, n2684, n2685, n2686, n2687, n2688, n2689, 
      n2690, n2691, n2692, n2693, n2694, n2695, n2696, n2697, n2698, n2699, 
      n2700, n2701, n2702, n2703, n2898, n2916, n2918, n2919, n2920, n2921, 
      n2996, n3029, n3030, n3033, n3035, n3038, n3040, n3043, n3045, n3048, 
      n3050, n3053, n3055, n3058, n3060, n3063, n3065, n3068, n3070, n3073, 
      n3075, n3078, n3080, n3083, n3085, n3088, n3090, n3093, n3095, n3098, 
      n3100, n3103, n3105, n3106, n3107, n3108, n3109, n3112, n3114, n3117, 
      n3121, n3125, n3129, n3133, n3137, n3141, n3145, n3149, n3153, n3157, 
      n3161, n3165, n3169, n3173, n3177, n3179, n3182, n3186, n3190, n3194, 
      n3198, n3202, n3206, n3210, n3214, n3218, n3222, n3226, n3230, n3234, 
      n3238, n3242, n3244, n3247, n3251, n3255, n3259, n3263, n3267, n3271, 
      n3275, n3279, n3283, n3287, n3291, n3295, n3299, n3303, n3307, n3309, 
      n3312, n3316, n3320, n3324, n3328, n3332, n3336, n3340, n3342, n3343, 
      n3346, n3348, n3351, n3353, n3356, n3358, n3359, n3362, n3364, n3367, 
      n3371, n3375, n3377, n3380, n3382, n3383, n3386, n3390, n3394, n3398, 
      n3400, n3403, n3405, n3406, n3409, n3413, n3415, n3416, n3417, n3418, 
      n3419, n3420, n3421, n3422, n3423, n3424, n3425, n3426, n3427, n3428, 
      n3429, n3430, n3431, n3432, n3433, n3434, n3435, n3436, n3437, n3438, 
      n3439, n3440, n3441, n3442, n3443, n3444, n3445, n3446, n3447, n3448, 
      n3449, n3450, n3451, n3452, n3453, n3454, n3455, n3456, n3457, n3458, 
      n3459, n3460, n3461, n3462, n3463, n3464, n3465, n3466, n3467, n3468, 
      n3469, n3470, n3471, n3472, n3473, n3474, n3475, n3476, n3477, n3478, 
      n3479, n3480, n3481, n3482, n3483, n3484, n3485, n3486, n3487, n3488, 
      n3489, n3490, n3491, n3492, n3493, n3494, n3495, n3496, n3497, n3498, 
      n3499, n3500, n3501, n3502, n3503, n3504, n3505, n3506, n3507, n3508, 
      n3509, n3510, n3511, n3512, n3513, n3514, n3515, n3516, n3517, n3518, 
      n3519, n3520, n3521, n3522, n3523, n3524, n3525, n3526, n3527, n3528, 
      n3529, n3530, n3531, n3532, n3533, n3534, n3535, n3536, n3537, n3538, 
      n3539, n3540, n3541, n3542, n3543, n3544, n3545, n3546, n3547, n3548, 
      n3549, n3550, n3551, n3552, n3553, n3554, n3555, n3556, n3557, n3558, 
      n3559, n3560, n3561, n3562, n3563, n3564, n3565, n3566, n3567, n3568, 
      n3569, n3570, n3571, n3572, n3573, n3574, n3575, n3576, n3577, n3578, 
      n3579, n3580, n3581, n3582, n3583, n3584, n3585, n3586, n3587, n3588, 
      n3589, n3590, n3591, n3592, n3593, n3594, n3595, n3596, n3597, n3598, 
      n3599, n3600, n3601, n3602, n3603, n3604, n3605, n3606, n3607, n3608, 
      n3609, n3610, n3611, n3612, n3613, n3614, n3615, n3616, n3617, n3618, 
      n3619, n3620, n3621, n3622, n3623, n3624, n3625, n3626, n3627, n3628, 
      n3629, n3630, n3631, n3632, n3633, n3634, n3635, n3636, n3637, n3638, 
      n3639, n3640, n3641, n3642, n3643, n3644, n3645, n3646, n3647, n3648, 
      n3649, n3650, n3651, n3652, n3653, n3654, n3655, n3656, n3657, n3658, 
      n3659, n3660, n3661, n3662, n3663, n3664, n3665, n3666, n3667, n3668, 
      n3669, n3670, n3671, n3672, n3673, n3674, n3675, n3676, n3677, n3678, 
      n3679, n3680, n3681, n3682, n3683, n3684, n3685, n3686, n3687, n3688, 
      n3689, n3690, n3691, n3692, n3693, n3694, n3695, n3696, n3697, n3698, 
      n3699, n3700, n3701, n3702, n3703, n3704, n3705, n3706, n3707, n3708, 
      n3709, n3710, n3711, n3712, n3713, n3714, n3715, n3716, n3717, n3718, 
      n3719, n3720, n3721, n3722, n3723, n3724, n3725, n3726, n3727, n3728, 
      n3729, n3730, n3731, n3732, n3733, n3734, n3735, n3736, n3737, n3738, 
      n3739, n3740, n3741, n3742, n3743, n3744, n3745, n3746, n3747, n3748, 
      n3749, n3750, n3751, n3752, n3753, n3754, n3755, n3756, n3757, n3758, 
      n3759, n3760, n3761, n3762, n3763, n3764, n3765, n3766, n3767, n3768, 
      n3769, n3770, n3771, n3772, n3773, n3774, n3775, n3776, n3777, n3778, 
      n3779, n3780, n3781, n3782, n3783, n3784, n3785, n3786, n3787, n3788, 
      n3789, n3790, n3791, n3792, n3793, n3794, n3795, n3796, n3797, n3798, 
      n3799, n3800, n3801, n3802, n3803, n3804, n3805, n3806, n3807, n3808, 
      n3809, n3810, n3811, n3812, n3813, n3814, n3815, n3816, n3817, n3818, 
      n3819, n3820, n3821, n3822, n3823, n3824, n3825, n3826, n3827, n3828, 
      n3829, n3830, n3831, n3832, n3833, n3834, n3835, n3836, n3837, n3838, 
      n3839, n3840, n3841, n3842, n3843, n3844, n3845, n3846, n3847, n3848, 
      n3849, n3850, n3851, n3852, n3853, n3854, n3855, n3856, n3857, n3858, 
      n3859, n3860, n3861, n3862, n3863, n3864, n3865, n3866, n3867, n3868, 
      n3869, n3870, n3871, n3872, n3873, n3874, n3875, n3876, n3877, n3878, 
      n3879, n3880, n3881, n3882, n3883, n3884, n3885, n3886, n3887, n3888, 
      n3889, n3890, n3891, n3892, n3893, n3894, n3895, n3896, n3897, n3898, 
      n3899, n3900, n3901, n3902, n3903, n3904, n3905, n3906, n3907, n3908, 
      n3909, n3910, n3911, n3912, n3913, n3914, n3915, n3916, n3917, n3918, 
      n3919, n3920, n3921, n3922, n3923, n3924, n3925, n3926, n3927, n3928, 
      n3929, n3930, n3931, n3932, n3933, n3934, n3935, n3936, n3937, n3938, 
      n3939, n3940, n3941, n3942, n3943, n3944, n3945, n3946, n3947, n3948, 
      n3949, n3950, n3951, n3952, n3953, n3954, n3955, n3956, n3957, n3958, 
      n3959, n3960, n3961, n3962, n3963, n3964, n3965, n3966, n3967, n3968, 
      n3969, n3970, n3971, n3972, n3973, n3974, n3975, n3976, n3977, n3978, 
      n3979, n3980, n3981, n3982, n3983, n3984, n3985, n3986, n3987, n3988, 
      n3989, n3990, n3991, n3992, n3993, n3994, n3995, n3996, n3997, n3998, 
      n3999, n4000, n4001, n4002, n4003, n4004, n4005, n4006, n4007, n4008, 
      n4009, n4010, n4011, n4012, n4013, n4014, n4015, n4016, n4017, n4018, 
      n4019, n4020, n4021, n4022, n4023, n4024, n4025, n4026, n4027, n4028, 
      n4029, n4030, n4031, n4032, n4033, n4034, n4035, n4036, n4037, n4038, 
      n4039, n4040, n4041, n4042, n4043, n4044, n4045, n4046, n4047, n4048, 
      n4049, n4050, n4051, n4052, n4053, n4054, n4055, n4056, n4057, n4058, 
      n4059, n4060, n4061, n4062, n4063, n4064, n4065, n4066, n4067, n4068, 
      n4069, n4070, n4071, n4072, n4073, n4074, n4075, n4076, n4077, n4078, 
      n4079, n4080, n4081, n4082, n4083, n4084, n4085, n4086, n4087, n4088, 
      n4089, n4090, n4091, n4092, n4093, n4094, n4095, n4096, n4097, n4098, 
      n4099, n4100, n4101, n4102, n4103, n4104, n4105, n4106, n4107, n4108, 
      n4109, n4110, n4111, n4112, n4113, n4114, n4115, n4116, n4117, n4118, 
      n4119, n4120, n4121, n4122, n4123, n4124, n4125, n4126, n4127, n4128, 
      n4129, n4130, n4131, n4132, n4133, n4134, n4135, n4136, n4137, n4138, 
      n4139, n4140, n4141, n4142, n4143, n4144, n4145, n4146, n4147, n4148, 
      n4149, n4150, n4151, n4152, n4153, n4154, n4155, n4156, n4157, n4158, 
      n4159, n4160, n4161, n4162, n4163, n4164, n4165, n4166, n4167, n4168, 
      n4169, n4170, n4171, n4172, n4173, n4174, n4175, n4176, n4177, n4178, 
      n4179, n4180, n4181, n4182, n4183, n4184, n4185, n4186, n4187, n4188, 
      n4189, n4190, n4191, n4192, n4193, n4194, n4195, n4196, n4197, n4198, 
      n4199, n4200, n4201, n4202, n4203, n4204, n4205, n4206, n4207, n4208, 
      n4209, n4210, n4211, n4212, n4213, n4214, n4215, n4216, n4217, n4218, 
      n4219, n4220, n4221, n4222, n4223, n4224, n4225, n4226, n4227, n4228, 
      n4229, n4230, n4231, n4232, n4233, n4234, n4235, n4236, n4237, n4238, 
      n4239, n4240, n4241, n4242, n4243, n4244, n4245, n4246, n4247, n4248, 
      n4249, n4250, n4251, n4252, n4253, n4254, n4255, n4256, n4257, n4258, 
      n4259, n4260, n4261, n4262, n4263, n4264, n4265, n4266, n4267, n4268, 
      n4269, n4270, n4271, n4272, n4273, n4274, n4275, n4276, n4277, n4278, 
      n4279, n4280, n4281, n4282, n4283, n4284, n4285, n4286, n4287, n4288, 
      n4289, n4290, n4291, n4292, n4293, n4294, n4295, n4296, n4297, n4298, 
      n4299, n4300, n4301, n4302, n4303, n4304, n4305, n4306, n4307, n4308, 
      n4309, n4310, n4311, n4312, n4313, n4314, n4315, n4316, n4317, n4318, 
      n4319, n4320, n4321, n4322, n4323, n4324, n4325, n4326, n4327, n4328, 
      n4329, n4330, n4331, n4332, n4333, n4334, n4335, n4336, n4337, n4338, 
      n4339, n4340, n4341, n4342, n4343, n4344, n4345, n4346, n4347, n4348, 
      n4349, n4350, n4351, n4352, n4353, n4354, n4355, n4356, n4357, n4358, 
      n4359, n4360, n4361, n4362, n4363, n4364, n4365, n4366, n4367, n4368, 
      n4369, n4370, n4371, n4372, n4373, n4374, n4375, n4376, n4377, n4378, 
      n4379, n4380, n4381, n4382, n4383, n4384, n4385, n4386, n4387, n4388, 
      n4389, n4390, n4391, n4392, n4393, n4394, n4395, n4396, n4397, n4398, 
      n4399, n4400, n4401, n4402, n4403, n4404, n4405, n4406, n4407, n4408, 
      n4409, n4410, n4411, n4412, n4413, n4414, n4415, n4416, n4417, n4418, 
      n4419, n4420, n4421, n4422, n4423, n4424, n4425, n4426, n4427, n4428, 
      n4429, n4430, n4431, n4432, n4433, n4434, n4435, n4436, n4437, n4438, 
      n4439, n4440, n4441, n4442, n4443, n4444, n4445, n4446, n4447, n4448, 
      n4449, n4450, n4451, n4452, n4453, n4454, n4455, n4456, n4457, n4458, 
      n4459, n4460, n4461, n4462, n4463, n4464, n4465, n4466, n4467, n4468, 
      n4469, n4470, n4471, n4472, n4473, n4474, n4475, n4476, n4477, n4478, 
      n4479, n4480, n4481, n4482, n4483, n4484, n4485, n4486, n4487, n4488, 
      n4489, n4490, n4491, n4492, n4493, n4494, n4495, n4496, n4497, n4498, 
      n4499, n4500, n4501, n4502, n4503, n4504, n4505, n4506, n4507, n4508, 
      n4509, n4510, n4511, n4512, n4513, n4514, n4515, n4516, n4517, n4518, 
      n4519, n4520, n4521, n4522, n4523, n4524, n4525, n4526, n4527, n4528, 
      n4529, n4530, n4531, n4532, n4533, n4534, n4535, n4536, n4537, n4538, 
      n4539, n4540, n4541, n4542, n4543, n4544, n4545, n4546, n4547, n4548, 
      n4549, n4550, n4551, n4552, n4553, n4554, n4555, n4556, n4557, n4558, 
      n4559, n4560, n4561, n4562, n4563, n4564, n4565, n4566, n4567, n4568, 
      n4569, n4570, n4571, n4572, n4573, n4574, n4575, n4576, n4577, n4578, 
      n4579, n4580, n4581, n4582, n4583, n4584, n4585, n4586, n4587, n4588, 
      n4589, n4590, n4591, n4592, n4593, n4594, n4595, n4596, n4597, n4598, 
      n4599, n4600, n4601, n4602, n4603, n4604, n4605, n4606, n4607, n4608, 
      n4609, n4610, n4611, n4612, n4613, n4614, n4615, n4616, n4617, n4618, 
      n4619, n4620, n4621, n4622, n4623, n4624, n4625, n4626, n4627, n4628, 
      n4629, n4630, n4631, n4632, n4633, n4634, n4635, n4636, n4637, n4638, 
      n4639, n4640, n4641, n4642, n4643, n4644, n4645, n4646, n4647, n4648, 
      n4649, n4650, n4651, n4652, n4653, n4654, n4655, n4656, n4657, n4658, 
      n4659, n4660, n4661, n4662, n4663, n4664, n4665, n4666, n4667, n4668, 
      n4669, n4670, n4671, n4672, n4673, n4674, n4675, n4676, n4677, n4678, 
      n4679, n4680, n4681, n4682, n4683, n4684, n4685, n4686, n4687, n4688, 
      n4689, n4690, n4691, n4692, n4693, n4694, n4695, n4696, n4697, n4698, 
      n4699, n4700, n4701, n4702, n4703, n4704, n4705, n4706, n4707, n4708, 
      n4709, n4710, n4711, n4712, n4713, n4714, n4715, n4716, n4717, n4718, 
      n4719, n4720, n4721, n4722, n4723, n4724, n4725, n4726, n4727, n4728, 
      n4729, n4730, n4731, n4732, n4733, n4734, n4735, n4736, n4737, n4738, 
      n4739, n4740, n4741, n4742, n4743, n4744, n4745, n4746, n4747, n4748, 
      n4749, n4750, n4751, n4752, n4753, n4754, n4755, n4756, n4757, n4758, 
      n4759, n4760, n4761, n4762, n4763, n4764, n4765, n4766, n4767, n4768, 
      n4769, n4770, n4771, n4772, n4773, n4774, n4775, n4776, n4777, n4778, 
      n4779, n4780, n4781, n4782, n4783, n4784, n4785, n4786, n4787, n4788, 
      n4789, n4790, n4791, n4792, n4793, n4794, n4795, n4796, n4797, n4798, 
      n4799, n4800, n4801, n4802, n4803, n4804, n4805, n4806, n4807, n4808, 
      n4809, n4810, n4811, n4812, n4813, n4814, n4815, n4816, n4817, n4818, 
      n4819, n4820, n4821, n4822, n4823, n4824, n4825, n4826, n4827, n4828, 
      n4829, n4830, n4831, n4832, n4833, n4834, n4835, n4836, n4837, n4838, 
      n4839, n4840, n4841, n4842, n4843, n4844, n4845, n4846, n4847, n4848, 
      n4849, n4850, n4851, n4852, n4853, n4854, n4855, n4856, n4857, n4858, 
      n4859, n4860, n4861, n4862, n4863, n4864, n4865, n4866, n4867, n4868, 
      n4869, n4870, n4871, n4872, n4873, n4874, n4875, n4876, n4877, n4878, 
      n4879, n4880, n4881, n4882, n4883, n4884, n4885, n4886, n4887, n4888, 
      n4889, n4890, n4891, n4892, n4893, n4894, n4895, n4896, n4897, n4898, 
      n4899, n4900, n4901, n4902, n4903, n4904, n4905, n4906, n4907, n4908, 
      n4909, n4910, n4911, n4912, n4913, n4914, n4915, n4916, n4917, n4918, 
      n4919, n4920, n4921, n4922, n4923, n4924, n4925, n4926, n4927, n4928, 
      n4929, n4930, n4931, n4932, n4933, n4934, n4935, n4936, n4937, n4938, 
      n4939, n4940, n4941, n4942, n4943, n4944, n4945, n4946, n4947, n4948, 
      n4949, n4950, n4951, n4952, n4953, n4954, n4955, n4956, n4957, n4958, 
      n4959, n4960, n4961, n4962, n4963, n4964, n4965, n4966, n4967, n4968, 
      n4969, n4970, n4971, n4972, n4973, n4974, n4975, n4976, n4977, n4978, 
      n4979, n4980, n4981, n4982, n4983, n4984, n4985, n4986, n4987, n4988, 
      n4989, n4990, n4991, n4992, n4993, n4994, n4995, n4996, n4997, n4998, 
      n4999, n5000, n5001, n5002, n5003, n5004, n5005, n5006, n5007, n5008, 
      n5009, n5010, n5011, n5012, n5013, n5014, n5015, n5016, n5017, n5018, 
      n5019, n5020, n5021, n5022, n5023, n5024, n5025, n5026, n5027, n5028, 
      n5029, n5030, n5031, n5032, n5033, n5034, n5035, n5036, n5037, n5038, 
      n5039, n5040, n5041, n5042, n5043, n5044, n5045, n5046, n5047, n5048, 
      n5049, n5050, n5051, n5052, n5053, n5054, n5055, n5056, n5057, n5058, 
      n5059, n5060, n5061, n5062, n5063, n5064, n5065, n5066, n5067, n5068, 
      n5069, n5070, n5071, n5072, n5073, n5074, n5075, n5076, n5077, n5078, 
      n5079, n5080, n5081, n5082, n5083, n5084, n5085, n5086, n5087, n5088, 
      n5089, n5090, n5091, n5092, n5093, n5094, n5095, n5096, n5097, n5098, 
      n5099, n5100, n5101, n5102, n5103, n5104, n5105, n5106, n5107, n5108, 
      n5109, n5110, n5111, n5112, n5113, n5114, n5115, n5116, n5117, n5118, 
      n5119, n5120, n5121, n5122, n5123, n5124, n5125, n5126, n5127, n5128, 
      n5129, n5130, n5131, n5132, n5133, n5134, n5135, n5136, n5137, n5138, 
      n5139, n5140, n5141, n5142, n5143, n5144, n5145, n5146, n5147, n5148, 
      n5149, n5150, n5151, n5152, n5153, n5154, n5155, n5156, n5157, n5158, 
      n5159, n5160, n5161, n5162, n5163, n5164, n5165, n5166, n5167, n5168, 
      n5169, n5170, n5171, n5172, n5173, n5174, n5175, n5176, n5177, n5178, 
      n5179, n5180, n5181, n5182, n5183, n5184, n5185, n5186, n5187, n5188, 
      n5189, n5190, n5191, n5192, n5193, n5194, n5195, n5196, n5197, n5198, 
      n5199, n5200, n5201, n5202, n5203, n5204, n5205, n5206, n5207, n5208, 
      n5209, n5210, n5211, n5212, n5213, n5214, n5215, n5216, n5217, n5218, 
      n5219, n5220, n5221, n5222, n5223, n5224, n5225, n5226, n5227, n5228, 
      n5229, n5230, n5231, n5232, n5233, n5234, n5235, n5236, n5237, n5238, 
      n5239, n5240, n5241, n5242, n5243, n5244, n5245, n5246, n5247, n5248, 
      n5249, n5250, n5251, n5252, n5253, n5254, n5255, n5256, n5257, n5258, 
      n5259, n5260, n5261, n5262, n5263, n5264, n5265, n5266, n5267, n5268, 
      n5269, n5270, n5271, n5272, n5273, n5274, n5275, n5276, n5277, n5278, 
      n5279, n5280, n5281, n5282, n5283, n5284, n5285, n5286, n5287, n5288, 
      n5289, n5290, n5291, n5292, n5293, n5294, n5295, n5296, n5297, n5298, 
      n5299, n5300, n5301, n5302, n5303, n5304, n5305, n5306, n5307, n5308, 
      n5309, n5310, n5311, n5312, n5313, n5314, n5315, n5316, n5317, n5318, 
      n5319, n5320, n5321, n5322, n5323, n5324, n5325, n5326, n5327, n5328, 
      n5329, n5330, n5331, n5332, n5333, n5334, n5335, n5336, n5337, n5338, 
      n5339, n5340, n5341, n5342, n5343, n5344, n5345, n5346, n5347, n5348, 
      n5349, n5350, n5351, n5352, n5353, n5354, n5355, n5356, n5357, n5358, 
      n5359, n5360, n5361, n5362, n5363, n5364, n5365, n5366, n5367, n5368, 
      n5369, n5370, n5371, n5372, n5373, n5374, n5375, n5376, n5377, n5378, 
      n5379, n5380, n5381, n5382, n5383, n5384, n5385, n5386, n5387, n5388, 
      n5389, n5390, n5391, n5392, n5393, n5394, n5395, n5396, n5397, n5398, 
      n5399, n5400, n5401, n5402, n5403, n5404, n5405, n5406, n5407, n5408, 
      n5409, n5410, n5411, n5412, n5413, n5414, n5415, n5416, n5417, n5418, 
      n5419, n5420, n5421, n5422, n5423, n5424, n5425, n5426, n5427, n5428, 
      n5429, n5430, n5431, n5432, n5433, n5434, n5435, n5436, n5437, n5438, 
      n5439, n5440, n5441, n5442, n5443, n5444, n5445, n5446, n5447, n5448, 
      n5449, n5450, n5451, n5452, n5453, n5454, n5455, n5456, n5457, n5458, 
      n5459, n5460, n5461, n5462, n5463, n5464, n5465, n5466, n5467, n5468, 
      n5469, n5470, n5471, n5472, n5473, n5474, n5475, n5476, n5477, n5478, 
      n5479, n5480, n5481, n5482, n5483, n5484, n5485, n5486, n5487, n5488, 
      n5489, n5490, n5491, n5492, n5493, n5494, n5495, n5496, n5497, n5498, 
      n5499, n5500, n5501, n5502, n5503, n5504, n5505, n5506, n5507, n5508, 
      n5509, n5510, n5511, n5512, n5513, n5514, n5515, n5516, n5517, n5518, 
      n5519, n5520, n5521, n5522, n5523, n5524, n5525, n5526, n5527, n5528, 
      n5529, n5530, n5531, n5532, n5533, n5534, n5535, n5536, n5537, n5538, 
      n5539, n5540, n5541, n5542, n5543, n5544, n5545, n5546, n5547, n5548, 
      n5549, n5550, n5551, n5552, n5553, n5554, n5555, n5556, n5557, n5558, 
      n5559, n5560, n5561, n5562, n5563, n5564, n5565, n5566, n5567, n5568, 
      n5569, n5570, n5571, n5572, n5573, n5574, n5575, n5576, n5577, n5578, 
      n5579, n5580, n5581, n5582, n5583, n5584, n5585, n5586, n5587, n5588, 
      n5589, n5590, n5591, n5592, n5593, n5594, n5595, n5596, n5597, n5598, 
      n5599, n5600, n5601, n5602, n5603, n5604, n5605, n5606, n5607, n5608, 
      n5609, n5610, n5611, n5612, n5613, n5614, n5615, n5616, n5617, n5618, 
      n5619, n5620, n5621, n5622, n5623, n5624, n5625, n5626, n5627, n5628, 
      n5629, n5630, n5631, n5632, n5633, n5634, n5635, n5636, n5637, n5638, 
      n5639, n5640, n5641, n5642, n5643, n5644, n5645, n5646, n5647, n5648, 
      n5649, n5650, n5651, n5652, n5653, n5654, n5655, n5656, n5657, n5658, 
      n5659, n5660, n5661, n5662, n5663, n5664, n5665, n5666, n5667, n5668, 
      n5669, n5670, n5671, n5672, n5673, n5674, n5675, n5676, n5677, n5678, 
      n5679, n5680, n5681, n5682, n5683, n5684, n5685, n5686, n5687, n5688, 
      n5689, n5690, n5691, n5692, n5693, n5694, n5695, n5696, n5697, n5698, 
      n5699, n5700, n5701, n5702, n5703, n5704, n5705, n5706, n5707, n5708, 
      n5709, n5710, n5711, n5712, n5713, n5714, n5715, n5716, n5717, n5718, 
      n5719, n5720, n5721, n5722, n5723, n5724, n5725, n5726, n5727, n5728, 
      n5729, n5730, n5731, n5732, n5733, n5734, n5735, n5736, n5737, n5738, 
      n5739, n5740, n5741, n5742, n5743, n5744, n5745, n5746, n5747, n5748, 
      n5749, n5750, n5751, n5752, n5753, n5754, n5755, n5756, n5757, n5758, 
      n5759, n5760, n5761, n5762, n5763, n5764, n5765, n5766, n5767, n5768, 
      n5769, n5770, n5771, n5772, n5773, n5774, n5775, n5776, n5777, n5778, 
      n5779, n5780, n5781, n5782, n5783, n5784, n5785, n5786, n5787, n5788, 
      n5789, n5790, n5791, n5792, n5793, n5794, n5795, n5796, n5797, n5798, 
      n5799, n5800, n5801, n5802, n5803, n5804, n5805, n5806, n5807, n5808, 
      n5809, n5810, n5811, n5812, n5813, n5814, n5815, n5816, n5817, n5818, 
      n5819, n5820, n5821, n5822, n5823, n5824, n5825, n5826, n5827, n5828, 
      n5829, n5830, n5831, n5832, n5833, n5834, n5835, n5836, n5837, n5838, 
      n5839, n5840, n5841, n5842, n5843, n5844, n5845, n5846, n5847, n5848, 
      n5849, n5850, n5851, n5852, n5853, n5854, n5855, n5856, n5857, n5858, 
      n5859, n5860, n5861, n5862, n5863, n5864, n5865, n5866, n5867, n5868, 
      n5869, n5870, n5871, n5872, n5873, n5874, n5875, n5876, n5877, n5878, 
      n5879, n5880, n5881, n5882, n5883, n5884, n5885, n5886, n5887, n5888, 
      n5889, n5890, n5891, n5892, n5893, n5894, n5895, n5896, n5897, n5898, 
      n5899, n5900, n5901, n5902, n5903, n5904, n5905, n5906, n5907, n5908, 
      n5909, n5910, n5911, n5912, n5913, n5914, n5915, n5916, n5917, n5918, 
      n5919, n5920, n5921, n5922, n5923, n5924, n5925, n5926, n5927, n5928, 
      n5929, n5930, n5931, n5932, n5933, n5934, n5935, n5936, n5937, n5938, 
      n5939, n5940, n5941, n5942, n5943, n5944, n5945, n5946, n5947, n5948, 
      n5949, n5950, n5951, n5952, n5953, n5954, n5955, n5956, n5957, n5958, 
      n5959, n5960, n5961, n5962, n5963, n5964, n5965, n5966, n5967, n5968, 
      n5969, n5970, n5971, n5972, n5973, n5974, n5975, n5976, n5977, n5978, 
      n5979, n5980, n5981, n5982, n5983, n5984, n5985, n5986, n5987, n5988, 
      n5989, n5990, n5991, n5992, n5993, n5994, n5995, n5996, n5997, n5998, 
      n5999, n6000, n6001, n6002, n6003, n6004, n6005, n6006, n6007, n6008, 
      n6009, n6010, n6011, n6012, n6013, n6014, n6015, n6016, n6017, n6018, 
      n6019, n6020, n6021, n6022, n6023, n6024, n6025, n6026, n6027, n6028, 
      n6029, n6030, n6031, n6032, n6033, n6034, n6035, n6036, n6037, n6038, 
      n6039, n6040, n6041, n6042, n6043, n6044, n6045, n6046, n6047, n6048, 
      n6049, n6050, n6051, n6052, n6053, n6054, n6055, n6056, n6057, n6058, 
      n6059, n6060, n6061, n6062, n6063, n6064, n6065, n6066, n6067, n6068, 
      n6069, n6070, n6071, n6072, n6073, n6074, n6075, n6076, n6077, n6078, 
      n6079, n6080, n6081, n6082, n6083, n6084, n6085, n6086, n6087, n6088, 
      n6089, n6090, n6091, n6092, n6093, n6094, n6095, n6096, n6097, n6098, 
      n6099, n6100, n6101, n6102, n6103, n6104, n6105, n6106, n6107, n6108, 
      n6109, n6110, n6111, n6112, n6113, n6114, n6115, n6116, n6117, n6118, 
      n6119, n6120, n6121, n6122, n6123, n6124, n6125, n6126, n6127, n6128, 
      n6129, n6130, n6131, n6132, n6133, n6134, n6135, n6136, n6137, n6138, 
      n6139, n6140, n6141, n6142, n6143, n6144, n6145, n6146, n6147, n6148, 
      n6149, n6150, n6151, n6152, n6153, n6154, n6155, n6156, n6157, n6158, 
      n6159, n6160, n6161, n6162, n6163, n6164, n6165, n6166, n6167, n6168, 
      n6169, n6170, n6171, n6172, n6173, n6174, n6175, n6176, n6177, n6178, 
      n6179, n6180, n6181, n6182, n6183, n6184, n6185, n6186, n6187, n6188, 
      n6189, n6190, n6191, n6192, n6193, n6194, n6195, n6196, n6197, n6198, 
      n6199, n6200, n6201, n6202, n6203, n6204, n6205, n6206, n6207, n6208, 
      n6209, n6210, n6211, n6212, n6213, n6214, n6215, n6216, n6217, n6218, 
      n6219, n6220, n6221, n6222, n6223, n6224, n6225, n6226, n6227, n6228, 
      n6229, n6230, n6231, n6232, n6233, n6234, n6235, n6236, n6237, n6238, 
      n6239, n6240, n6241, n6242, n6243, n6244, n6245, n6246, n6247, n6248, 
      n6249, n6250, n6251, n6252, n6253, n6254, n6255, n6256, n6257, n6258, 
      n6259, n6260, n6261, n6262, n6263, n6264, n6265, n6266, n6267, n6268, 
      n6269, n6270, n6271, n6272, n6273, n6274, n6275, n6276, n6277, n6278, 
      n6279, n6280, n6281, n6282, n6283, n6284, n6285, n6286, n6287, n6288, 
      n6289, n6290, n6291, n6292, n6293, n6294, n6295, n6296, n6297, n6298, 
      n6299, n6300, n6301, n6302, n6303, n6304, n6305, n6306, n6307, n6308, 
      n6309, n6310, n6311, n6312, n6313, n6314, n6315, n6316, n6317, n6318, 
      n6319, n6320, n6321, n6322, n6323, n6324, n6325, n6326, n6327, n6328, 
      n6329, n6330, n6331, n6332, n6333, n6334, n6335, n6336, n6337, n6338, 
      n6339, n6340, n6341, n6342, n6343, n6344, n6345, n6346, n6347, n6348, 
      n6349, n6350, n6351, n6352, n6353, n6354, n6355, n6356, n6357, n6358, 
      n6359, n6360, n6361, n6362, n6363, n6364, n6365, n6366, n6367, n6368, 
      n6369, n6370, n6371, n6372, n6373, n6374, n6375, n6376, n6377, n6378, 
      n6379, n6380, n6381, n6382, n6383, n6384, n6385, n6386, n6387, n6388, 
      n6389, n6390, n6391, n6392, n6393, n6394, n6395, n6396, n6397, n6398, 
      n6399, n6400, n6401, n6402, n6403, n6404, n6405, n6406, n6407, n6408, 
      n6409, n6410, n6411, n6412, n6413, n6414, n6415, n6416, n6417, n6418, 
      n6419, n6420, n6421, n6422, n6423, n6424, n6425, n6426, n6427, n6428, 
      n6429, n6430, n6431, n6432, n6433, n6434, n6435, n6436, n6437, n6438, 
      n6439, n6440, n6441, n6442, n6443, n6444, n6445, n6446, n6447, n6448, 
      n6449, n6450, n6451, n6452, n6453, n6454, n6455, n6456, n6457, n6458, 
      n6459, n6460, n6461, n6462, n6463, n6464, n6465, n6466, n6467, n6468, 
      n6469, n6470, n6471, n6472, n6473, n6474, n6475, n6476, n6477, n6478, 
      n6479, n6480, n6481, n6482, n6483, n6484, n6485, n6486, n6487, n6488, 
      n6489, n6490, n6491, n6492, n6493, n6494, n6495, n6496, n6497, n6498, 
      n6499, n6500, n6501, n6502, n6503, n6504, n6505, n6506, n6507, n6508, 
      n6509, n6510, n6511, n6512, n6513, n6514, n6515, n6516, n6517, n6518, 
      n6519, n6520, n6521, n6522, n6523, n6524, n6525, n6526, n6527, n6528, 
      n6529, n6530, n6531, n6532, n6533, n6534, n6535, n6536, n6537, n6538, 
      n6539, n6540, n6541, n6542, n6543, n6544, n6545, n6546, n6547, n6548, 
      n6549, n6550, n6551, n6552, n6553, n6554, n6555, n6556, n6557, n6558, 
      n6559, n6560, n6561, n6562, n6563, n6564, n6565, n6566, n6567, n6568, 
      n6569, n6570, n6571, n6572, n6573, n6574, n6575, n6576, n6577, n6578, 
      n6579, n6580, n6581, n6582, n6583, n6584, n6585, n6586, n6587, n6588, 
      n6589, n6590, n6591, n6592, n6593, n6594, n6595, n6596, n6597, n6598, 
      n6599, n6600, n6601, n6602, n6603, n6604, n6605, n6606, n6607, n6608, 
      n6609, n6610, n6611, n6612, n6613, n6614, n6615, n6616, n6617, n6618, 
      n6619, n6620, n6621, n6622, n6623, n6624, n6625, n6626, n6627, n6628, 
      n6629, n6630, n6631, n6632, n6633, n6634, n6635, n6636, n6637, n6638, 
      n6639, n6640, n6641, n6642, n6643, n6644, n6645, n6646, n6647, n6648, 
      n6649, n6650, n6651, n6652, n6653, n6654, n6655, n6656, n6657, n6658, 
      n6659, n6660, n6661, n6662, n6663, n6664, n6665, n6666, n6667, n6668, 
      n6669, n6670, n6671, n6672, n6673, n6674, n6675, n6676, n6677, n6678, 
      n6679, n6680, n6681, n6682, n6683, n6684, n6685, n6686, n6687, n6688, 
      n6689, n6690, n6691, n6692, n6693, n6694, n6695, n6696, n6697, n6698, 
      n6699, n6700, n6701, n6702, n6703, n6704, n6705, n6706, n6707, n6708, 
      n6709, n6710, n6711, n6712, n6713, n6714, n6715, n6716, n6717, n6718, 
      n6719, n6720, n6721, n6722, n6723, n6724, n6725, n6726, n6727, n6728, 
      n6729, n6730, n6731, n6732, n6733, n6734, n6735, n6736, n6737, n6738, 
      n6739, n6740, n6741, n6742, n6743, n6744, n6745, n6746, n6747, n6748, 
      n6749, n6750, n6751, n6752, n6753, n6754, n6755, n6756, n6757, n6758, 
      n6759, n6760, n6761, n6762, n6763, n6764, n6765, n6766, n6767, n6768, 
      n6769, n6770, n6771, n6772, n6773, n6774, n6775, n6776, n6777, n6778, 
      n6779, n6780, n6781, n6782, n6783, n6784, n6785, n6786, n6787, n6788, 
      n6789, n6790, n6791, n6792, n6793, n6794, n6795, n6796, n6797, n6798, 
      n6799, n6800, n6801, n6802, n6803, n6804, n6805, n6806, n6807, n6808, 
      n6809, n6810, n6811, n6812, n6813, n6814, n6815, n6816, n6817, n6818, 
      n6819, n6820, n6821, n6822, n6823, n6824, n6825, n6826, n6827, n6828, 
      n6829, n6830, n6831, n6832, n6833, n6834, n6835, n6836, n6837, n6838, 
      n6839, n6840, n6841, n6842, n6843, n6844, n6845, n6846, n6847, n6848, 
      n6849, n6850, n6851, n6852, n6853, n6854, n6855, n6856, n6857, n6858, 
      n6859, n6860, n6861, n6862, n6863, n6864, n6865, n6866, n6867, n6868, 
      n6869, n6870, n6871, n6872, n6873, n6874, n6875, n6876, n6877, n6878, 
      n6879, n6880, n6881, n6882, n6883, n6884, n6885, n6886, n6887, n6888, 
      n6889, n6890, n6891, n6892, n6893, n6894, n6895, n6896, n6897, n6898, 
      n6899, n6900, n6901, n6902, n6903, n6904, n6905, n6906, n6907, n6908, 
      n6909, n6910, n6911, n6912, n6913, n6914, n6915, n6916, n6917, n6918, 
      n6919, n6920, n6921, n6922, n6923, n6924, n6925, n6926, n6927, n6928, 
      n6929, n6930, n6931, n6932, n6933, n6934, n6935, n6936, n6937, n6938, 
      n6939, n6940, n6941, n6942, n6943, n6944, n6945, n6946, n6947, n6948, 
      n6949, n6950, n6951, n6952, n6953, n6954, n6955, n6956, n6957, n6958, 
      n6959, n6960, n6961, n6962, n6963, n6964, n6965, n6966, n6967, n6968, 
      n6969, n6970, n6971, n6972, n6973, n6974, n6975, n6976, n6977, n6978, 
      n6979, n6980, n6981, n6982, n6983, n6984, n6985, n6986, n6987, n6988, 
      n6989, n6990, n6991, n6992, n6993, n6994, n6995, n6996, n6997, n6998, 
      n6999, n7000, n7001, n7002, n7003, n7004, n7005, n7006, n7007, n7008, 
      n7009, n7010, n7011, n7012, n7013, n7014, n7015, n7016, n7017, n7018, 
      n7019, n7020, n7021, n7022, n7023, n7024, n7025, n7026, n7027, n7028, 
      n7029, n7030, n7031, n7032, n7033, n7034, n7035, n7036, n7037, n7038, 
      n7039, n7040, n7041, n7042, n7043, n7044, n7045, n7046, n7047, n7048, 
      n7049, n7050, n7051, n7052, n7053, n7054, n7055, n7056, n7057, n7058, 
      n7059, n7060, n7061, n7062, n7063, n7064, n7065, n7066, n7067, n7068, 
      n7069, n7070, n7071, n7072, n7073, n7074, n7075, n7076, n7077, n7078, 
      n7079, n7080, n7081, n7082, n7083, n7084, n7085, n7086, n7087, n7088, 
      n7089, n7090, n7091, n7092, n7093, n7094, n7095, n7096, n7097, n7098, 
      n7099, n7100, n7101, n7102, n7103, n7104, n7105, n7106, n7107, n7108, 
      n7109, n7110, n7111, n7112, n7113, n7114, n7115, n7116, n7117, n7118, 
      n7119, n7120, n7121, n7122, n7123, n7124, n7125, n7126, n7127, n7128, 
      n7129, n7130, n7131, n7132, n7133, n7134, n7135, n7136, n7137, n7138, 
      n7139, n7140, n7141, n7142, n7143, n7144, n7145, n7146, n7147, n7148, 
      n7149, n7150, n7151, n7152, n7153, n7154, n7155, n7156, n7157, n7158, 
      n7159, n7160, n7161, n7162, n7163, n7164, n7165, n7166, n7167, n7168, 
      n7169, n7170, n7171, n7172, n7173, n7174, n7175, n7176, n7177, n7178, 
      n7179, n7180, n7181, n7182, n7183, n7184, n7185, n7186, n7187, n7188, 
      n7189, n7190, n7191, n7192, n7193, n7194, n7195, n7196, n7197, n7198, 
      n7199, n7200, n7201, n7202, n7203, n7204, n7205, n7206, n7207, n7208, 
      n7209, n7210, n7211, n7212, n7213, n7214, n7215, n7216, n7217, n7218, 
      n7219, n7220, n7221, n7222, n7223, n7224, n7225, n7226, n7227, n7228, 
      n7229, n7230, n7231, n7232, n7233, n7234, n7235, n7236, n7237, n7238, 
      n7239, n7240, n7241, n7242, n7243, n7244, n7245, n7246, n7247, n7248, 
      n7249, n7250, n7251, n7252, n7253, n7254, n7255, n7256, n7257, n7258, 
      n7259, n7260, n7261, n7262, n7263, n7264, n7265, n7266, n7267, n7268, 
      n7269, n7270, n7271, n7272, n7273, n7274, n7275, n7276, n7277, n7278, 
      n7279, n7280, n7281, n7282, n7283, n7284, n7285, n7286, n7287, n7288, 
      n7289, n7290, n7291, n7292, n7293, n7294, n7295, n7296, n7297, n7298, 
      n7299, n7300, n7301, n7302, n7303, n7304, n7305, n7306, n7307, n7308, 
      n7309, n7310, n7311, n7312, n7313, n7314, n7315, n7316, n7317, n7318, 
      n7319, n7320, n7321, n7322, n7323, n7324, n7325, n7326, n7327, n7328, 
      n7329, n7330, n7331, n7332, n7333, n7334, n7335, n7336, n7337, n7338, 
      n7339, n7340, n7341, n7342, n7343, n7344, n7345, n7346, n7347, n7348, 
      n7349, n7350, n7351, n7352, n7353, n7354, n7355, n7356, n7357, n7358, 
      n7359, n7360, n7361, n7362, n7363, n7364, n7365, n7366, n7367, n7368, 
      n7369, n7370, n7371, n7372, n7373, n7374, n7375, n7376, n7377, n7378, 
      n7379, n7380, n7381, n7382, n7383, n7384, n7385, n7386, n7387, n7388, 
      n7389, n7390, n7391, n7392, n7393, n7394, n7395, n7396, n7397, n7398, 
      n7399, n7400, n7401, n7402, n7403, n7404, n7405, n7406, n7407, n7408, 
      n7409, n7410, n7411, n7412, n7413, n7414, n7415, n7416, n7417, n7418, 
      n7419, n7420, n7421, n7422, n7423, n7424, n7425, n7426, n7427, n7428, 
      n7429, n7430, n7431, n7432, n7433, n7434, n7435, n7436, n7437, n7438, 
      n7439, n7440, n7441, n7442, n7443, n7444, n7445, n7446, n7447, n7448, 
      n7449, n7450, n7451, n7452, n7453, n7454, n7455, n7456, n7457, n7458, 
      n7459, n7460, n7461, n7462, n7463, n7464, n7465, n7466, n7467, n7468, 
      n7469, n7470, n7471, n7472, n7473, n7474, n7475, n7476, n7477, n7478, 
      n7479, n7480, n7481, n7482, n7483, n7484, n7485, n7486, n7487, n7488, 
      n7489, n7490, n7491, n7492, n7493, n7494, n7495, n7496, n7497, n7498, 
      n7499, n7500, n7501, n7502, n7503, n7504, n7505, n7506, n7507, n7508, 
      n7509, n7510, n7511, n7512, n7513, n7514, n7515, n7516, n7517, n7518, 
      n7519, n7520, n7521, n7522, n7523, n7524, n7525, n7526, n7527, n7528, 
      n7529, n7530, n7531, n7532, n7533, n7534, n7535, n7536, n7537, n7538, 
      n7539, n7540, n7541, n7542, n7543, n7544, n7545, n7546, n7547, n7548, 
      n7549, n7550, n7551, n7552, n7553, n7554, n7555, n7556, n7557, n7558, 
      n7559, n7560, n7561, n7562, n7563, n7564, n7565, n7566, n7567, n7568, 
      n7569, n7570, n7571, n7572, n7573, n7574, n7575, n7576, n7577, n7578, 
      n7579, n7580, n7581, n7582, n7583, n7584, n7585, n7586, n7587, n7588, 
      n7589, n7590, n7591, n7592, n7593, n7594, n7595, n7596, n7597, n7598, 
      n7599, n7600, n7601, n7602, n7603, n7604, n7605, n7606, n7607, n7608, 
      n7609, n7610, n7611, n7612, n7613, n7614, n7615, n7616, n7617, n7618, 
      n7619, n7620, n7621, n7622, n7623, n7624, n7625, n7626, n7627, n7628, 
      n7629, n7630, n7631, n7632, n7633, n7634, n7635, n7636, n7637, n7638, 
      n7639, n7640, n7641, n7642, n7643, n7644, n7645, n7646, n7647, n7648, 
      n7649, n7650, n7651, n7652, n7653, n7654, n7655, n7656, n7657, n7658, 
      n7659, n7660, n7661, n7662, n7663, n7664, n7665, n7666, n7667, n7668, 
      n7669, n7670, n7671, n7672, n7673, n7674, n7675, n7676, n7677, n7678, 
      n7679, n7680, n7681, n7682, n7683, n7684, n7685, n7686, n7687, n7688, 
      n7689, n7690, n7691, n7692, n7693, n7694, n7695, n7696, n7697, n7698, 
      n7699, n7700, n7701, n7702, n7703, n7704, n7705, n7706, n7707, n7708, 
      n7709, n7710, n7711, n7712, n7713, n7714, n7715, n7716, n7717, n7718, 
      n7719, n7720, n7721, n7722, n7723, n7724, n7725, n7726, n7727, n7728, 
      n7729, n7730, n7731, n7732, n7733, n7734, n7735, n7736, n7737, n7738, 
      n7739, n7740, n7741, n7742, n7743, n7744, n7745, n7746, n7747, n7748, 
      n7749, n7750, n7751, n7752, n7753, n7754, n7755, n7756, n7757, n7758, 
      n7759, n7760, n7761, n7762, n7763, n7764, n7765, n7766, n7767, n7768, 
      n7769, n7770, n7771, n7772, n7773, n7774, n7775, n7776, n7777, n7778, 
      n7779, n7780, n7781, n7782, n7783, n7784, n7785, n7786, n7787, n7788, 
      n7789, n7790, n7791, n7792, n7793, n7794, n7795, n7796, n7797, n7798, 
      n7799, n7800, n7801, n7802, n7803, n7804, n7805, n7806, n7807, n7808, 
      n7809, n7810, n7811, n7812, n7813, n7814, n7815, n7816, n7817, n7818, 
      n7819, n7820, n7821, n7822, n7823, n7824, n7825, n7826, n7827, n7828, 
      n7829, n7830, n7831, n7832, n7833, n7834, n7835, n7836, n7837, n7838, 
      n7839, n7840, n7841, n7842, n7843, n7844, n7845, n7846, n7847, n7848, 
      n7849, n7850, n7851, n7852, n7853, n7854, n7855, n7856, n7857, n7858, 
      n7859, n7860, n7861, n7862, n7863, n7864, n7865, n7866, n7867, n7868, 
      n7869, n7870, n7871, n7872, n7873, n7874, n7875, n7876, n7877, n7878, 
      n7879, n7880, n7881, n7882, n7883, n7884, n7885, n7886, n7887, n7888, 
      n7889, n7890, n7891, n7892, n7893, n7894, n7895, n7896, n7897, n7898, 
      n7899, n7900, n7901, n7902, n7903, n7904, n7905, n7906, n7907, n7908, 
      n7909, n7910, n7911, n7912, n7913, n7914, n7915, n7916, n7917, n7918, 
      n7919, n7920, n7921, n7922, n7923, n7924, n7925, n7926, n7927, n7928, 
      n7929, n7930, n7931, n7932, n7933, n7934, n7935, n7936, n7937, n7938, 
      n7939, n7940, n7941, n7942, n7943, n7944, n7945, n7946, n7947, n7948, 
      n7949, n7950, n7951, n7952, n7953, n7954, n7955, n7956, n7957, n7958, 
      n7959, n7960, n7961, n7962, n7963, n7964, n7965, n7966, n7967, n7968, 
      n7969, n7970, n7971, n7972, n7973, n7974, n7975, n7976, n7977, n7978, 
      n7979, n7980, n7981, n7982, n7983, n7984, n7985, n7986, n7987, n7988, 
      n7989, n7990, n7991, n7992, n7993, n7994, n7995, n7996, n7997, n7998, 
      n7999, n8000, n8001, n8002, n8003, n8004, n8005, n8006, n8007, n8008, 
      n8009, n8010, n8011, n8012, n8013, n8014, n8015, n8016, n8017, n8018, 
      n8019, n8020, n8021, n8022, n8023, n8024, n8025, n8026, n8027, n8028, 
      n8029, n8030, n8031, n8032, n8033, n8034, n8035, n8036, n8037, n8038, 
      n8039, n8040, n8041, n8042, n8043, n8044, n8045, n8046, n8047, n8048, 
      n8049, n8050, n8051, n8052, n8053, n8054, n8055, n8056, n8057, n8058, 
      n8059, n8060, n8061, n8062, n8063, n8064, n8065, n8066, n8067, n8068, 
      n8069, n8070, n8071, n8072, n8073, n8074, n8075, n8076, n8077, n8078, 
      n8079, n8080, n8081, n8082, n8083, n8084, n8085, n8086, n8087, n8088, 
      n8089, n8090, n8091, n8092, n8093, n8094, n8095, n8096, n8097, n8098, 
      n8099, n8100, n8101, n8102, n8103, n8104, n8105, n8106, n8107, n8108, 
      n8109, n8110, n8111, n8112, n8113, n8114, n8115, n8116, n8117, n8118, 
      n8119, n8120, n8121, n8122, n8123, n8124, n8125, n8126, n8127, n8128, 
      n8129, n8130, n8131, n8132, n8133, n8134, n8135, n8136, n8137, n8138, 
      n8139, n8140, n8141, n8142, n8143, n8144, n8145, n8146, n8147, n8148, 
      n8149, n8150, n8151, n8152, n8153, n8154, n8155, n8156, n8157, n8158, 
      n8159, n8160, n8161, n8162, n8163, n8164, n8165, n8166, n8167, n8168, 
      n8169, n8170, n8171, n8172, n8173, n8174, n8175, n8176, n8177, n8178, 
      n8179, n8180, n8181, n8182, n8183, n8184, n8185, n8186, n8187, n8188, 
      n8189, n8190, n8191, n8192, n8193, n8194, n8195, n8196, n8197, n8198, 
      n8199, n8200, n8201, n8202, n8203, n8204, n8205, n8206, n8207, n8208, 
      n8209, n8210, n8211, n8212, n8213, n8214, n8215, n8216, n8217, n8218, 
      n8219, n8220, n8221, n8222, n8223, n8224, n8225, n8226, n8227, n8228, 
      n8229, n8230, n8231, n8232, n8233, n8234, n8235, n8236, n8237, n8238, 
      n8239, n8240, n8241, n8242, n8243, n8244, n8245, n8246, n8247, n8248, 
      n8249, n8250, n8251, n8252, n8253, n8254, n8255, n8256, n8257, n8258, 
      n8259, n8260, n8261, n8262, n8263, n8264, n8265, n8266, n8267, n8268, 
      n8269, n8270, n8271, n8272, n8273, n8274, n8275, n8276, n8277, n8278, 
      n8279, n8280, n8281, n8282, n8283, n8284, n8285, n8286, n8287, n8288, 
      n8289, n8290, n8291, n8292, n8293, n8294, n8295, n8296, n8297, n8298, 
      n8299, n8300, n8301, n8302, n8303, n8304, n8305, n8306, n8307, n8308, 
      n8309, n8310, n8311, n8312, n8313, n8314, n8315, n8316, n8317, n8318, 
      n8319, n8320, n8321, n8322, n8323, n8324, n8325, n8326, n8327, n8328, 
      n8329, n8330, n8331, n8332, n8333, n8334, n8335, n8336, n8337, n8338, 
      n8339, n8340, n8341, n8342, n8343, n8344, n8345, n8346, n8347, n8348, 
      n8349, n8350, n8351, n8352, n8353, n8354, n8355, n8356, n8357, n8358, 
      n8359, n8360, n8361, n8362, n8363, n8364, n8365, n8366, n8367, n8368, 
      n8369, n8370, n8371, n8372, n8373, n8374, n8375, n8376, n8377, n8378, 
      n8379, n8380, n8381, n8382, n8383, n8384, n8385, n8386, n8387, n8388, 
      n8389, n8390, n8391, n8392, n8393, n8394, n8395, n8396, n8397, n8398, 
      n8399, n8400, n8401, n8402, n8403, n8404, n8405, n8406, n8407, n8408, 
      n8409, n8410, n8411, n8412, n8413, n8414, n8415_port, n8416, n8417_port, 
      n8418_port, n8419_port, n8420_port, n8421_port, n8422_port, n8423_port, 
      n8424, n8425, n8426, n8427_port, n8428_port, n8429_port, n8430_port, 
      n8431, n8432, n8433, n8434, n8435, n8436, n8437, n8438, n8439, n8440, 
      n8441, n8442, n8443, n8444, n8445, n8446, n8447, n8448, n8449, n8450, 
      n8451, n8452, n8453, n8454, n8455, n8456, n8457, n8458, n8459, n8460, 
      n8461, n8462, n8463, n8464, n8465, n8466, n8467, n8468, n8469, n8470, 
      n8471, n8472, n8473, n8474, n8475, n8476, n8477, n8478, n8479, n8480, 
      n8481, n8482, n8483, n8484, n8485, n8486, n8487, n8488, n8489, n8490, 
      n8491, n8492, n8493, n8494, n8495, n8496, n8497, n8498, n8499, n8500, 
      n8501, n8502, n8503, n8504, n8505, n8506, n8507, n8508, n8509, n8510, 
      n8511, n8512, n8513, n8514, n8515, n8516, n8517, n8518, n8519, n8520, 
      n8521, n8522, n8523, n8524, n8525, n8526, n8527, n8528, n8529, n8530, 
      n8531, n8532, n8533, n8534, n8535, n8536, n8537, n8538, n8539, n8540, 
      n8541, n8542, n8543, n8544, n8545, n8546, n8547, n8548, n8549, n8550, 
      n8551, n8552, n8553, n8554, n8555, n8556, n8557, n8558, n8559_port, n8560
      , n8561_port, n8562_port, n8563_port, n8564_port, n8565_port, n8566_port,
      n8567_port, n8568, n8569, n8570, n8571_port, n8572_port, n8573_port, 
      n8574_port, n8575, n8576, n8577, n8578, n8579, n8580, n8581, n8582, n8583
      , n8584, n8585, n8586, n8587, n8588, n8589, n8590, n8591, n8592, n8593, 
      n8594, n8595, n8596, n8597, n8598, n8599, n8600, n8601, n8602, n8603, 
      n8604, n8605, n8606, n8607, n8608, n8609, n8610, n8611, n8612, n8613, 
      n8614, n8615, n8616, n8617, n8618, n8619, n8620, n8621, n8622, n8623, 
      n8624, n8625, n8626, n8627, n8628, n8629, n8630, n8631, n8632, n8633, 
      n8634, n8635, n8636, n8637, n8638, n8639, n8640, n8641, n8642, n8643, 
      n8644, n8645, n8646, n8647, n8648, n8649, n8650, n8651, n8652, n8653, 
      n8654, n8655, n8656, n8657, n8658, n8659, n8660, n8661, n8662, n8663, 
      n8664, n8665, n8666, n8667, n8668, n8669, n8670, n8671, n8672, n8673, 
      n8674, n8675, n8676, n8677, n8678, n8679, n8680, n8681, n8682, n8683, 
      n8684, n8685, n8686, n8687, n8688, n8689, n8690, n8691, n8692, n8693, 
      n8694, n8695, n8696, n8697, n8698, n8699, n8700, n8701, n8702_port, 
      n8703_port, n8704_port, n8705_port, n8706_port, n8707_port, n8708_port, 
      n8709_port, n8710_port, n8711_port, n8712_port, n8713_port, n8714_port, 
      n8715_port, n8716_port, n8717_port, n8718_port, n8719_port, n8720_port, 
      n8721_port, n8722_port, n8723_port, n8724_port, n8725_port, n8726_port, 
      n8727_port, n8728_port, n8729_port, n8730_port, n8731_port, n8732_port, 
      n8733_port, n8734_port, n8735_port, n8736_port, n8737_port, n8738_port, 
      n8739_port, n8740_port, n8741_port, n8742_port, n8743_port, n8744_port, 
      n8745_port, n8746_port, n8747_port, n8748_port, n8749_port, n8750_port, 
      n8751_port, n8752_port, n8753_port, n8754_port, n8755_port, n8756_port, 
      n8757_port, n8758_port, n8759_port, n8760_port, n8761_port, n8762_port, 
      n8763_port, n8764_port, n8765_port, n8766_port, n8767_port, n8768, n8769,
      n8770, n8771, n8772, n8773, n8774, n8775, n8776, n8777, n8778, n8779, 
      n8780, n8781, n8782, n8783, n8784, n8785, n8786, n8787_port, n8788_port, 
      n8789_port, n8790_port, n8791_port, n8792, n8793, n8794, n8795, n8796, 
      n8797, n8798, n8799, n8800, n8801, n8802, n8803, n8804, n8805, n8806, 
      n8807, n8808, n8809, n8810, n8811, n8812, n8813, n8814, n8815, n8816, 
      n8817, n8818, n8819, n8820, n8821, n8822, n8823, n8824, n8825, n8826, 
      n8827, n8828, n8829, n8830, n8831, n8832, n8833_port, n8834_port, n8835, 
      n8836, n8837, n8838, n8839, n8840, n8841, n8842, n8843, n8844, n8845, 
      n8846, n8847, n8848, n8849, n8850, n8851, n8852, n8853, n8854, n8855, 
      n8856, n8857, n8858, n8859, n8860, n8861, n8862, n8863, n8864, n8865, 
      n8866, n8867, n8868, n8869, n8870, n8871, n8872, n8873, n8874, n8875, 
      n8876, n8877, n8878, n8879, n8880, n8881, n8882, n8883, n8884, n8885, 
      n8886, n8887, n8888, n8889, n8890, n8891, n8892, n8893, n8894, n8895, 
      n8896, n8897, n8898, n8899, n8900, n8901, n8902, n8903, n8904, n8905, 
      n8906, n8907, n8908, n8909, n8910, n8911, n8912, n8913, n8914, n8915, 
      n8916, n8917, n8918, n8919, n8920, n8921, n8922, n8923, n8924, n8925, 
      n8926, n8927, n8928, n8929, n8930, n8931, n8932, n8933, n8934, n8935, 
      n8936, n8937, n8938, n8939, n8940, n8941, n8942, n8943, n8944, n8945, 
      n8946, n8947, n8948, n8949, n8950, n8951, n8952, n8953, n8954, n8955, 
      n8956, n8957, n8958, n8959, n8960, n8961, n8962, n8963, n8964, n8965, 
      n8966, n8967, n8968, n8969, n8970, n8971, n8972, n8973, n8974, n8975, 
      n8976, n8977, n8978, n8979, n8980, n8981, n8982, n8983, n8984, n8985, 
      n8986, n8987, n8988, n8989, n8990, n8991, n8992, n8993, n8994, n8995, 
      n8996, n8997, n8998, n8999, n9000, n9001, n9002, n9003, n9004, n9005, 
      n9006, n9007, n9008, n9009, n9010, n9011, n9012, n9013, n9014, n9015, 
      n9016, n9017, n9018, n9019, n9020, n9021, n9022, n9023, n9024, n9025, 
      n9026, n9027, n9028, n9029, n9030, n9031, n9032, n9033, n9034, n9035, 
      n9036, n9037, n9038, n9039, n9040, n9041, n9042, n9043, n9044, n9045, 
      n9046, n9047, n9048, n9049, n9050, n9051, n9052, n9053, n9054, n9055, 
      n9056, n9057, n9058, n9059, n9060, n9061, n9062, n9063, n9064, n9065, 
      n9066, n9067, n9068, n9069, n9070, n9071, n9072, n9073, n9074, n9075, 
      n9076, n9077, n9078, n9079, n9080, n9081, n9082, n9083, n9084, n9085, 
      n9086, n9087, n9088, n9089, n9090, n9091, n9092, n9093, n9094, n9095, 
      n9096, n9097, n9098, n9099, n9100, n9101, n9102, n9103, n9104, n9105, 
      n9106, n9107, n9108, n9109, n9110, n9111, n9112, n9113, n9114, n9115, 
      n9116, n9117, n9118, n9119, n9120, n9121, n9122, n9123, n9124, n9125, 
      n9126, n9127, n9128, n9129, n9130, n9131, n9132, n9133, n9134, n9135, 
      n9136, n9137, n9138, n9139, sub_189_carry_6_port, n1, n2, n3, n4, n5, n6,
      n8, n9, n10, n12, n13, n14, n15, n16, n18, n19, n20, n21, n22, n23, n24, 
      n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39
      , n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, 
      n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68
      , n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n432, n433, n434
      , n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446,
      n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, n458, 
      n459, n460, n461, n462, n463, n464, n465, n466, n467, n468, n469, n470, 
      n471, n472, n473, n474, n475, n476, n477, n478, n479, n480, n481, n482, 
      n483, n484, n485, n486, n487, n488, n489, n490, n491, n492, n493, n494, 
      n495, n592, n593, n594, n595, n596, n597, n598, n599, n600, n601, n602, 
      n603, n604, n605, n606, n607, n608, n609, n610, n611, n612, n613, n614, 
      n615, n616, n617, n618, n619, n620, n621, n622, n623, n624, n625, n626, 
      n627, n628, n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, 
      n639, n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, 
      n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662, 
      n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673, n674, 
      n675, n676, n677, n678, n679, n680, n681, n682, n683, n684, n685, n686, 
      n687, n688, n689, n690, n691, n692, n693, n694, n695, n696, n697, n698, 
      n699, n700, n701, n702, n703, n704, n705, n706, n707, n708, n709, n710, 
      n711, n712, n713, n714, n715, n716, n717, n718, n719, n720, n721, n722, 
      n723, n724, n725, n726, n727, n728, n729, n730, n731, n732, n733, n734, 
      n735, n736, n737, n738, n739, n740, n741, n742, n743, n744, n745, n746, 
      n747, n748, n749, n750, n751, n752, n753, n754, n755, n756, n757, n758, 
      n759, n760, n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, 
      n771, n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782, 
      n783, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144, 
      n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154, 
      n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164, 
      n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174, 
      n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184, 
      n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194, 
      n1195, n1196, n1197, n1198, n1199, n1296, n1297, n1298, n1299, n1300, 
      n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, 
      n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, 
      n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, 
      n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, 
      n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, 
      n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, 
      n1361, n1362, n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, 
      n1371, n1372, n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380, 
      n1381, n1382, n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390, 
      n1391, n1392, n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400, 
      n1401, n1402, n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410, 
      n1411, n1412, n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420, 
      n1421, n1422, n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430, 
      n1431, n1432, n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440, 
      n1441, n1442, n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450, 
      n1451, n1452, n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460, 
      n1461, n1462, n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470, 
      n1471, n1472, n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480, 
      n1481, n1482, n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490, 
      n1491, n1492, n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500, 
      n1501, n1502, n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510, 
      n1511, n1512, n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520, 
      n1521, n1522, n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530, 
      n1531, n1532, n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540, 
      n1541, n1542, n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550, 
      n1551, n1648, n1649, n1650, n1651, n1652, n1653, n1654, n1655, n1656, 
      n1657, n1658, n1659, n1660, n1661, n1662, n1663, n1664, n1665, n1666, 
      n1667, n1668, n1669, n1670, n1671, n1672, n1673, n1674, n1675, n1676, 
      n1677, n1678, n1679, n1680, n1681, n1682, n1683, n1684, n1685, n1686, 
      n1687, n1688, n1689, n1690, n1691, n1692, n1693, n1694, n1695, n1696, 
      n1697, n1698, n1699, n1700, n1701, n1702, n1703, n1704, n1705, n1706, 
      n1707, n1708, n1709, n1710, n1711, n1712, n1713, n1714, n1715, n1716, 
      n1717, n1718, n1719, n1720, n1721, n1722, n1723, n1724, n1725, n1726, 
      n1727, n1728, n1729, n1730, n1731, n1732, n1733, n1734, n1735, n1736, 
      n1737, n1738, n1739, n1740, n1741, n1742, n1743, n1744, n1745, n1746, 
      n1747, n1748, n1749, n1750, n1751, n1752, n1753, n1754, n1755, n1756, 
      n1757, n1758, n1759, n1760, n1761, n1762, n1763, n1764, n1765, n1766, 
      n1767, n1768, n1769, n1770, n1771, n1772, n1773, n1774, n1775, n1776, 
      n1777, n1778, n1779, n1780, n1781, n1782, n1783, n1784, n1785, n1786, 
      n1787, n1788, n1789, n1790, n1791, n1792, n1793, n1794, n1795, n1796, 
      n1797, n1798, n1799, n1800, n1801, n1802, n1803, n1804, n1805, n1806, 
      n1807, n1808, n1809, n1810, n1811, n1812, n1813, n1814, n1815, n1816, 
      n1817, n1818, n1819, n1820, n1821, n1822, n1823, n1824, n1825, n1826, 
      n1827, n1828, n1829, n1830, n1831, n1832, n1833, n1834, n1835, n1836, 
      n1837, n1838, n1839, n2544, n2545, n2546, n2547, n2548, n2549, n2550, 
      n2551, n2552, n2553, n2554, n2555, n2556, n2557, n2558, n2559, n2560, 
      n2561, n2562, n2563, n2564, n2565, n2566, n2567, n2568, n2569, n2570, 
      n2571, n2572, n2573, n2574, n2575, n2576, n2577, n2578, n2579, n2580, 
      n2581, n2582, n2583, n2584, n2585, n2586, n2587, n2588, n2589, n2590, 
      n2591, n2592, n2593, n2594, n2595, n2596, n2597, n2598, n2599, n2600, 
      n2601, n2602, n2603, n2604, n2605, n2606, n2607, n2704, n2705, n2706, 
      n2707, n2708, n2709, n2710, n2711, n2712, n2713, n2714, n2715, n2716, 
      n2717, n2718, n2719, n2720, n2721, n2722, n2723, n2724, n2725, n2726, 
      n2727, n2728, n2729, n2730, n2731, n2732, n2733, n2734, n2735, n2736, 
      n2737, n2738, n2739, n2740, n2741, n2742, n2743, n2744, n2745, n2746, 
      n2747, n2748, n2749, n2750, n2751, n2752, n2753, n2754, n2755, n2756, 
      n2757, n2758, n2759, n2760, n2761, n2762, n2763, n2764, n2765, n2766, 
      n2767, n2768, n2769, n2770, n2771, n2772, n2773, n2774, n2775, n2776, 
      n2777, n2778, n2779, n2780, n2781, n2782, n2783, n2784, n2785, n2786, 
      n2787, n2788, n2789, n2790, n2791, n2792, n2793, n2794, n2795, n2796, 
      n2797, n2798, n2799, n2800, n2801, n2802, n2803, n2804, n2805, n2806, 
      n2807, n2808, n2809, n2810, n2811, n2812, n2813, n2814, n2815, n2816, 
      n2817, n2818, n2819, n2820, n2821, n2822, n2823, n2824, n2825, n2826, 
      n2827, n2828, n2829, n2830, n2831, n2832, n2833, n2834, n2835, n2836, 
      n2837, n2838, n2839, n2840, n2841, n2842, n2843, n2844, n2845, n2846, 
      n2847, n2848, n2849, n2850, n2851, n2852, n2853, n2854, n2855, n2856, 
      n2857, n2858, n2859, n2860, n2861, n2862, n2863, n2864, n2865, n2866, 
      n2867, n2868, n2869, n2870, n2871, n2872, n2873, n2874, n2875, n2876, 
      n2877, n2878, n2879, n2880, n2881, n2882, n2883, n2884, n2885, n2886, 
      n2887, n2888, n2889, n2890, n2891, n2892, n2893, n2894, n2895, n2896, 
      n2897, n2899, n2900, n2901, n2902, n2903, n2904, n2905, n2906, n2907, 
      n2908, n2909, n2910, n2911, n2912, n2913, n2914, n2915, n2917, n2922, 
      n2923, n2924, n2925, n2926, n2927, n2928, n2929, n2930, n2931, n2932, 
      n2933, n2934, n2935, n2936, n2937, n2938, n2939, n2940, n2941, n2942, 
      n2943, n2944, n2945, n2946, n2947, n2948, n2949, n2950, n2951, n2952, 
      n2953, n2954, n2955, n2956, n2957, n2958, n2959, n2960, n2961, n2962, 
      n2963, n2964, n2965, n2966, n2967, n2968, n2969, n2970, n2971, n2972, 
      n2973, n2974, n2975, n2976, n2977, n2978, n2979, n2980, n2981, n2982, 
      n2983, n2984, n2985, n2986, n2987, n2988, n2989, n2990, n2991, n2992, 
      n2993, n2994, n2995, n2997, n2998, n2999, n3000, n3001, n3002, n3003, 
      n3004, n3005, n3006, n3007, n3008, n3009, n3010, n3011, n3012, n3013, 
      n3014, n3015, n3016, n3017, n3018, n3019, n3020, n3021, n3022, n3023, 
      n3024, n3025, n3026, n3027, n3028, n3031, n3032, n3034, n3036, n3037, 
      n3039, n3041, n3042, n3044, n3046, n3047, n3049, n3051, n3052, n3054, 
      n3056, n3057, n3059, n3061, n3062, n3064, n3066, n3067, n3069, n3071, 
      n3072, n3074, n3076, n3077, n3079, n3081, n3082, n3084, n3086, n3087, 
      n3089, n3091, n3092, n3094, n3096, n3097, n3099, n3101, n3102, n3104, 
      n3110, n3111, n3113, n3115, n3116, n3118, n3119, n3120, n3122, n3123, 
      n3124, n3126, n3127, n3128, n3130, n3131, n3132, n3134, n3135, n3136, 
      n3138, n3139, n3140, n3142, n3143, n3144, n3146, n3147, n3148, n3150, 
      n3151, n3152, n3154, n3155, n3156, n3158, n3159, n3160, n3162, n3163, 
      n3164, n3166, n3167, n3168, n3170, n3171, n3172, n3174, n3175, n3176, 
      n3178, n3180, n3181, n3183, n3184, n3185, n3187, n3188, n3189, n3191, 
      n3192, n3193, n3195, n3196, n3197, n3199, n3200, n3201, n3203, n3204, 
      n3205, n3207, n3208, n3209, n3211, n3212, n3213, n3215, n3216, n3217, 
      n3219, n3220, n3221, n3223, n3224, n3225, n3227, n3228, n3229, n3231, 
      n3232, n3233, n3235, n3236, n3237, n3239, n3240, n3241, n3243, n3245, 
      n3246, n3248, n3249, n3250, n3252, n3253, n3254, n3256, n3257, n3258, 
      n3260, n3261, n3262, n3264, n3265, n3266, n3268, n3269, n3270, n3272, 
      n3273, n3274, n3276, n3277, n3278, n3280, n3281, n3282, n3284, n3285, 
      n3286, n3288, n3289, n3290, n3292, n3293, n3294, n3296, n3297, n3298, 
      n3300, n3301, n3302, n3304, n3305, n3306, n3308, n3310, n3311, n3313, 
      n3314, n3315, n3317, n3318, n3319, n3321, n3322, n3323, n3325, n3326, 
      n3327, n3329, n3330, n3331, n3333, n3334, n3335, n3337, n3338, n3339, 
      n3341, n3344, n3345, n3347, n3349, n3350, n3352, n3354, n3355, n3357, 
      n3360, n3361, n3363, n3365, n3366, n3368, n3369, n3370, n3372, n3373, 
      n3374, n3376, n3378, n3379, n3381, n3384, n3385, n3387, n3388, n3389, 
      n3391, n3392, n3393, n3395, n3396, n3397, n3399, n3401, n3402, n3404, 
      n3407, n3408, n3410, n3411, n3412, n3414, n9140, n9141, n9142, n9143, 
      n9144, n9145, n9146, n9147, n9148, n9149, n9150, n9151, n9152, n9153, 
      n9154, n9155, n9156, n9157, n9158, n9159, n9160, n9161, n9162, n9163, 
      n9164, n9165, n9166, n9167, n9168, n9169, n9170, n9171, n9172, n9173, 
      n9174, n9175, n9176, n9177, n9178, n9179, n9180, n9181, n9182, n9183, 
      n9184, n9185, n9186, n9187, n9188, n9189, n9190, n9191, n9192, n9193, 
      n9194, n9195, n9196, n9197, n9198, n9199, n9200, n9201, n9202, n9203, 
      n9204, n9205, n9206, n9207, n9208, n9209, n9210, n9211, n9212, n9213, 
      n9214, n9215, n9216, n9217, n9218, n9219, n9220, n9221, n9222, n9223, 
      n9224, n9225, n9226, n9227, n9228, n9229, n9230, n9231, n9232, n9233, 
      n9234, n9235, n9236, n9237, n9238, n9239, n9240, n9241, n9242, n9243, 
      n9244, n9245, n9246, n9247, n9248, n9249, n9250, n9251, n9252, n9253, 
      n9254, n9255, n9256, n9257, n9258, n9259, n9260, n9261, n9262, n9263, 
      n9264, n9265, n9266, n9267, n9268, n9269, n9270, n9271, n9272, n9273, 
      n9274, n9275, n9276, n9277, n9278, n9279, n9280, n9281, n9282, n9283, 
      n9284, n9285, n9286, n9287, n9288, n9289, n9290, n9291, n9292, n9293, 
      n9294, n9295, n9296, n9297, n9298, n9299, n9300, n9301, n9302, n9303, 
      n9304, n9305, n9306, n9307, n9308, n9309, n9310, n9311, n9312, n9313, 
      n9314, n9315, n9316, n9317, n9318, n9319, n9320, n9321, n9322, n9323, 
      n9324, n9325, n9326, n9327, n9328, n9329, n9330, n9331, n9332, n9333, 
      n9334, n9335, n9336, n9337, n9338, n9339, n9340, n9341, n9342, n9343, 
      n9344, n9345, n9346, n9347, n9348, n9349, n9350, n9351, n9352, n9353, 
      n9354, n9355, n9356, n9357, n9358, n9359, n9360, n9361, n9362, n9363, 
      n9364, n9365, n9366, n9367, n9368, n9369, n9370, n9371, n9372, n9373, 
      n9374, n9375, n9376, n9377, n9378, n9379, n9380, n9381, n9382, n9383, 
      n9384, n9385, n9386, n9387, n9388, n9389, n9390, n9391, n9392, n9393, 
      n9394, n9395, n9396, n9397, n9398, n9399, n9400, n9401, n9402, n9403, 
      n9404, n9405, n9406, n9407, n9408, n9409, n9410, n9411, n9412, n9413, 
      n9414, n9415, n9416, n9417, n9418, n9419, n9420, n9421, n9422, n9423, 
      n9424, n9425, n9426, n9427, n9428, n9429, n9430, n9431, n9432, n9433, 
      n9434, n9435, n9436, n9437, n9438, n9439, n9440, n9441, n9442, n9443, 
      n9444, n9445, n9446, n9447, n9448, n9449, n9450, n9451, n9452, n9453, 
      n9454, n9455, n9456, n9457, n9458, n9459, n9460, n9461, n9462, n9463, 
      n9464, n9465, n9466, n9467, n9468, n9469, n9470, n9471, n9472, n9473, 
      n9474, n9475, n9476, n9477, n9478, n9479, n9480, n9481, n9482, n9483, 
      n9484, n9485, n9486, n9487, n9488, n9489, n9490, n9491, n9492, n9493, 
      n9494, n9495, n9496, n9497, n9498, n9499, n9500, n9501, n9502, n9503, 
      n9504, n9505, n9506, n9507, n9508, n9509, n9510, n9511, n9512, n9513, 
      n9514, n9515, n9516, n9517, n9518, n9519, n9520, n9521, n9522, n9523, 
      n9524, n9525, n9526, n9527, n9528, n9529, n9530, n9531, n9532, n9533, 
      n9534, n9535, n9536, n9537, n9538, n9539, n9540, n9541, n9542, n9543, 
      n9544, n9545, n9546, n9547, n9548, n9549, n9550, n9551, n9552, n9553, 
      n9554, n9555, n9556, n9557, n9558, n9559, n9560, n9561, n9562, n9563, 
      n9564, n9565, n9566, n9567, n9568, n9569, n9570, n9571, n9572, n9573, 
      n9574, n9575, n9576, n9577, n9578, n9579, n9580, n9581, n9582, n9583, 
      n9584, n9585, n9586, n9587, n9588, n9589, n9590, n9591, n9592, n9593, 
      n9594, n9595, n9596, n9597, n9598, n9599, n9600, n9601, n9602, n9603, 
      n9604, n9605, n9606, n9607, n9608, n9609, n9610, n9611, n9612, n9613, 
      n9614, n9615, n9616, n9617, n9618, n9619, n9620, n9621, n9622, n9623, 
      n9624, n9625, n9626, n9627, n9628, n9629, n9630, n9631, n9632, n9633, 
      n9634, n9635, n9636, n9637, n9638, n9639, n9640, n9641, n9642, n9643, 
      n9644, n9645, n9646, n9647, n9648, n9649, n9650, n9651, n9652, n9653, 
      n9654, n9655, n9656, n9657, n9658, n9659, n9660, n9661, n9662, n9663, 
      n9664, n9665, n9666, n9667, n9668, n9669, n9670, n9671, n9672, n9673, 
      n9674, n9675, n9676, n9677, n9678, n9679, n9680, n9681, n9682, n9683, 
      n9684, n9685, n9686, n9687, n9688, n9689, n9690, n9691, n9692, n9693, 
      n9694, n9695, n9696, n9697, n9698, n9699, n9700, n9701, n9702, n9703, 
      n9704, n9705, n9706, n9707, n9708, n9709, n9710, n9711, n9712, n9713, 
      n9714, n9715, n9716, n9717, n9718, n9719, n9720, n9721, n9722, n9723, 
      n9724, n9725, n9726, n9727, n9728, n9729, n9730, n9731, n9732, n9733, 
      n9734, n9735, n9736, n9737, n9738, n9739, n9740, n9741, n9742, n9743, 
      n9744, n9745, n9746, n9747, n9748, n9749, n9750, n9751, n9752, n9753, 
      n9754, n9755, n9756, n9757, n9758, n9759, n9760, n9761, n9762, n9763, 
      n9764, n9765, n9766, n9767, n9768, n9769, n9770, n9771, n9772, n9773, 
      n9774, n9775, n9776, n9777, n9778, n9779, n9780, n9781, n9782, n9783, 
      n9784, n9785, n9786, n9787, n9788, n9789, n9790, n9791, n9792, n9793, 
      n9794, n9795, n9796, n9797, n9798, n9799, n9800, n9801, n9802, n9803, 
      n9804, n9805, n9806, n9807, n9808, n9809, n9810, n9811, n9812, n9813, 
      n9814, n9815, n9816, n9817, n9818, n9819, n9820, n9821, n9822, n9823, 
      n9824, n9825, n9826, n9827, n9828, n9829, n9830, n9831, n9832, n9833, 
      n9834, n9835, n9836, n9837, n9838, n9839, n9840, n9841, n9842, n9843, 
      n9844, n9845, n9846, n9847, n9848, n9849, n9850, n9851, n9852, n9853, 
      n9854, n9855, n9856, n9857, n9858, n9859, n9860, n9861, n9862, n9863, 
      n9864, n9865, n9866, n9867, n9868, n9869, n9870, n9871, n9872, n9873, 
      n9874, n9875, n9876, n9877, n9878, n9879, n9880, n9881, n9882, n9883, 
      n9884, n9885, n9886, n9887, n9888, n9889, n9890, n9891, n9892, n9893, 
      n9894, n9895, n9896, n9897, n9898, n9899, n9900, n9901, n9902, n9903, 
      n9904, n9905, n9906, n9907, n9908, n9909, n9910, n9911, n9912, n9913, 
      n9914, n9915, n9916, n9917, n9918, n9919, n9920, n9921, n9922, n9923, 
      n9924, n9925, n9926, n9927, n9928, n9929, n9930, n9931, n9932, n9933, 
      n9934, n9935, n9936, n9937, n9938, n9939, n9940, n9941, n9942, n9943, 
      n9944, n9945, n9946, n9947, n9948, n9949, n9950, n9951, n9952, n9953, 
      n9954, n9955, n9956, n9957, n9958, n9959, n9960, n9961, n9962, n9963, 
      n9964, n9965, n9966, n9967, n9968, n9969, n9970, n9971, n9972, n9973, 
      n9974, n9975, n9976, n9977, n9978, n9979, n9980, n9981, n9982, n9983, 
      n9984, n9985, n9986, n9987, n9988, n9989, n9990, n9991, n9992, n9993, 
      n9994, n9995, n9996, n9997, n9998, n9999, n10000, n10001, n10002, n10003,
      n10004, n10005, n10006, n10007, n10008, n10009, n10010, n10011, n10012, 
      n10013, n10014, n10015, n10016, n10017, n10018, n10019, n10020, n10021, 
      n10022, n10023, n10024, n10025, n10026, n10027, n10028, n10029, n10030, 
      n10031, n10032, n10033, n10034, n10035, n10036, n10037, n10038, n10039, 
      n10040, n10041, n10042, n10043, n10044, n10045, n10046, n10047, n10048, 
      n10049, n10050, n10051, n10052, n10053, n10054, n10055, n10056, n10057, 
      n10058, n10059, n10060, n10061, n10062, n10063, n10064, n10065, n10066, 
      n10067, n10068, n10069, n10070, n10071, n10072, n10073, n10074, n10075, 
      n10076, n10077, n10078, n10079, n10080, n10081, n10082, n10083, n10084, 
      n10085, n10086, n10087, n10088, n10089, n10090, n10091, n10092, n10093, 
      n10094, n10095, n10096, n10097, n10098, n10099, n10100, n10101, n10102, 
      n10103, n10104, n10105, n10106, n10107, n10108, n10109, n10110, n10111, 
      n10112, n10113, n10114, n10115, n10116, n10117, n10118, n10119, n10120, 
      n10121, n10122, n10123, n10124, n10125, n10126, n10127, n10128, n10129, 
      n10130, n10131, n10132, n10133, n10134, n10135, n10136, n10137, n10138, 
      n10139, n10140, n10141, n10142, n10143, n10144, n10145, n10146, n10147, 
      n10148, n10149, n10150, n10151, n10152, n10153, n10154, n10155, n10156, 
      n10157, n10158, n10159, n10160, n10161, n10162, n10163, n10164, n10165, 
      n10166, n10167, n10168, n10169, n10170, n10171, n10172, n10173, n10174, 
      n10175, n10176, n10177, n10178, n10179, n10180, n10181, n10182, n10183, 
      n10184, n10185, n10186, n10187, n10188, n10189, n10190, n10191, n10192, 
      n10193, n10194, n10195, n10196, n10197, n10198, n10199, n10200, n10201, 
      n10202, n10203, n10204, n10205, n10206, n10207, n10208, n10209, n10210, 
      n10211, n10212, n10213, n10214, n10215, n10216, n10217, n10218, n10219, 
      n10220, n10221, n10222, n10223, n10224, n10225, n10226, n10227, n10228, 
      n10229, n10230, n10231, n10232, n10233, n10234, n10235, n10236, n10237, 
      n10238, n10239, n10240, n10241, n10242, n10243, n10244, n10245, n10246, 
      n10247, n10248, n10249, n10250, n10251, n10252, n10253, n10254, n10255, 
      n10256, n10257, n10258, n10259, n10260, n10261, n10262, n10263, n10264, 
      n10265, n10266, n10267, n10268, n10269, n10270, n10271, n10272, n10273, 
      n10274, n10275, n10276, n10277, n10278, n10279, n10280, n10281, n10282, 
      n10283, n10284, n10285, n10286, n10287, n10288, n10289, n10290, n10291, 
      n10292, n10293, n10294, n10295, n10296, n10297, n10298, n10299, n10300, 
      n10301, n10302, n10303, n10304, n10305, n10306, n10307, n10308, n10309, 
      n10310, n10311, n10312, n10313, n10314, n10315, n10316, n10317, n10318, 
      n10319, n10320, n10321, n10322, n10323, n10324, n10325, n10326, n10327, 
      n10328, n10329, n10330, n10331, n10332, n10333, n10334, n10335, n10336, 
      n10337, n10338, n10339, n10340, n10341, n10342, n10343, n10344, n10345, 
      n10346, n10347, n10348, n10349, n10350, n10351, n10352, n10353, n10354, 
      n10355, n10356, n10357, n10358, n10359, n10360, n10361, n10362, n10363, 
      n10364, n10365, n10366, n10367, n10368, n10369, n10370, n10371, n10372, 
      n10373, n10374, n10375, n10376, n10377, n10378, n10379, n10380, n10381, 
      n10382, n10383, n10384, n10385, n10386, n10387, n10388, n10389, n10390, 
      n10391, n10392, n10393, n10394, n10395, n10396, n10397, n10398, n10399, 
      n10400, n10401, n10402, n10403, n10404, n10405, n10406, n10407, n10408, 
      n10409, n10410, n10411, n10412, n10413, n10414, n10415, n10416, n10417, 
      n10418, n10419, n10420, n10421, n10422, n10423, n10424, n10425, n10426, 
      n10427, n10428, n10429, n10430, n10431, n10432, n10433, n10434, n10435, 
      n10436, n10437, n10438, n10439, n10440, n10441, n10442, n10443, n10444, 
      n10445, n10446, n10447, n10448, n10449, n10450, n10451, n10452, n10453, 
      n10454, n10455, n10456, n10457, n10458, n10459, n10460, n10461, n10462, 
      n10463, n10464, n10465, n10466, n10467, n10468, n10469, n10470, n10471, 
      n10472, n10473, n10474, n10475, n10476, n10477, n10478, n10479, n10480, 
      n10481, n10482, n10483, n10484, n10485, n10486, n10487, n10488, n10489, 
      n10490, n10491, n10492, n10493, n10494, n10495, n10496, n10497, n10498, 
      n10499, n10500, n10501, n10502, n10503, n10504, n10505, n10506, n10507, 
      n10508, n10509, n10510, n10511, n10512, n10513, n10514, n10515, n10516, 
      n10517, n10518, n10519, n10520, n10521, n10522, n10523, n10524, n10525, 
      n10526, n10527, n10528, n10529, n10530, n10531, n10532, n10533, n10534, 
      n10535, n10536, n10537, n10538, n10539, n10540, n10541, n10542, n10543, 
      n10544, n10545, n10546, n10547, n10548, n10549, n10550, n10551, n10552, 
      n10553, n10554, n10555, n10556, n10557, n10558, n10559, n10560, n10561, 
      n10562, n10563, n10564, n10565, n10566, n10567, n10568, n10569, n10570, 
      n10571, n10572, n10573, n10574, n10575, n10576, n10577, n10578, n10579, 
      n10580, n10581, n10582, n10583, n10584, n10585, n10586, n10587, n10588, 
      n10589, n10590, n10591, n10592, n10593, n10594, n10595, n10596, n10597, 
      n10598, n10599, n10600, n10601, n10602, n10603, n10604, n10605, n10606, 
      n10607, n10608, n10609, n10610, n10611, n10612, n10613, n10614, n10615, 
      n10616, n10617, n10618, n10619, n10620, n10621, n10622, n10623, n10624, 
      n10625, n10626, n10627, n10628, n10629, n10630, n10631, n10632, n10633, 
      n10634, n10635, n10636, n10637, n10638, n10639, n10640, n10641, n10642, 
      n10643, n10644, n10645, n10646, n10647, n10648, n10649, n10650, n10651, 
      n10652, n10653, n10654, n10655, n10656, n10657, n10658, n10659, n10660, 
      n10661, n10662, n10663, n10664, n10665, n10666, n10667, n10668, n10669, 
      n10670, n10671, n10672, n10673, n10674, n10675, n10676, n10677, n10678, 
      n10679, n10680, n10681, n10682, n10683, n10684, n10685, n10686, n10687, 
      n10688, n10689, n10690, n10691, n10692, n10693, n10694, n10695, n10696, 
      n10697, n10698, n10699, n10700, n10701, n10702, n10703, n10704, n10705, 
      n10706, n10707, n10708, n10709, n10710, n10711, n10712, n10713, n10714, 
      n10715, n10716, n10717, n10718, n10719, n10720, n10721, n10722, n10723, 
      n10724, n10725, n10726, n10727, n10728, n10729, n10730, n10731, n10732, 
      n10733, n10734, n10735, n10736, n10737, n10738, n10739, n10740, n10741, 
      n10742, n10743, n10744, n10745, n10746, n10747, n10748, n10749, n10750, 
      n10751, n10752, n10753, n10754, n10755, n10756, n10757, n10758, n10759, 
      n10760, n10761, n10762, n10763, n10764, n10765, n10766, n10767, n10768, 
      n10769, n10770, n10771, n10772, n10773, n10774, n10775, n10776, n10777, 
      n10778, n10779, n10780, n10781, n10782, n10783, n10784, n10785, n10786, 
      n10787, n10788, n10789, n10790, n10791, n10792, n10793, n10794, n10795, 
      n10796, n10797, n10798, n10799, n10800, n10801, n10802, n10803, n10804, 
      n10805, n10806, n10807, n10808, n10809, n10810, n10811, n10812, n10813, 
      n10814, n10815, n10816, n10817, n10818, n10819, n10820, n10821, n10822, 
      n10823, n10824, n10825, n10826, n10827, n10828, n10829, n10830, n10831, 
      n10832, n10833, n10834, n10835, n10836, n10837, n10838, n10839, n10840, 
      n10841, n10842, n10843, n10844, n10845, n10846, n10847, n10848, n10849, 
      n10850, n10851, n10852, n10853, n10854, n10855, n10856, n10857, n10858, 
      n10859, n10860, n10861, n10862, n10863, n10864, n10865, n10866, n10867, 
      n10868, n10869, n10870, n10871, n10872, n10873, n10874, n10875, n10876, 
      n10877, n10878, n10879, n10880, n10881, n10882, n10883, n10884, n10885, 
      n10886, n10887, n10888, n10889, n10890, n10891, n10892, n10893, n10894, 
      n10895, n10896, n10897, n10898, n10899, n10900, n10901, n10902, n10903, 
      n10904, n10905, n10906, n10907, n10908, n10909, n10910, n10911, n10912, 
      n10913, n10914, n10915, n10916, n10917, n10918, n10919, n10920, n10921, 
      n_1185, n_1186, n_1187, n_1188, n_1189, n_1190, n_1191, n_1192, n_1193, 
      n_1194, n_1195, n_1196, n_1197, n_1198, n_1199, n_1200, n_1201, n_1202, 
      n_1203, n_1204, n_1205, n_1206, n_1207, n_1208, n_1209, n_1210, n_1211, 
      n_1212, n_1213, n_1214, n_1215, n_1216, n_1217, n_1218, n_1219, n_1220, 
      n_1221, n_1222, n_1223, n_1224, n_1225, n_1226, n_1227, n_1228, n_1229, 
      n_1230, n_1231, n_1232, n_1233, n_1234, n_1235, n_1236, n_1237, n_1238, 
      n_1239, n_1240, n_1241, n_1242, n_1243, n_1244, n_1245, n_1246, n_1247, 
      n_1248, n_1249, n_1250, n_1251, n_1252, n_1253, n_1254, n_1255, n_1256, 
      n_1257, n_1258, n_1259, n_1260, n_1261, n_1262, n_1263, n_1264, n_1265, 
      n_1266, n_1267, n_1268, n_1269, n_1270, n_1271, n_1272, n_1273, n_1274, 
      n_1275, n_1276, n_1277, n_1278, n_1279, n_1280, n_1281, n_1282, n_1283, 
      n_1284, n_1285, n_1286, n_1287, n_1288, n_1289, n_1290, n_1291, n_1292, 
      n_1293, n_1294, n_1295, n_1296, n_1297, n_1298, n_1299, n_1300, n_1301, 
      n_1302, n_1303, n_1304, n_1305, n_1306, n_1307, n_1308, n_1309, n_1310, 
      n_1311, n_1312, n_1313, n_1314, n_1315, n_1316, n_1317, n_1318, n_1319, 
      n_1320, n_1321, n_1322, n_1323, n_1324, n_1325, n_1326, n_1327, n_1328, 
      n_1329, n_1330, n_1331, n_1332, n_1333, n_1334, n_1335, n_1336, n_1337, 
      n_1338, n_1339, n_1340, n_1341, n_1342, n_1343, n_1344, n_1345, n_1346, 
      n_1347, n_1348, n_1349, n_1350, n_1351, n_1352, n_1353, n_1354, n_1355, 
      n_1356, n_1357, n_1358, n_1359, n_1360, n_1361, n_1362, n_1363, n_1364, 
      n_1365, n_1366, n_1367, n_1368, n_1369, n_1370, n_1371, n_1372, n_1373, 
      n_1374, n_1375, n_1376, n_1377, n_1378, n_1379, n_1380, n_1381, n_1382, 
      n_1383, n_1384, n_1385, n_1386, n_1387, n_1388, n_1389, n_1390, n_1391, 
      n_1392, n_1393, n_1394, n_1395, n_1396, n_1397, n_1398, n_1399, n_1400, 
      n_1401, n_1402, n_1403, n_1404, n_1405, n_1406, n_1407, n_1408, n_1409, 
      n_1410, n_1411, n_1412, n_1413, n_1414, n_1415, n_1416, n_1417, n_1418, 
      n_1419, n_1420, n_1421, n_1422, n_1423, n_1424, n_1425, n_1426, n_1427, 
      n_1428, n_1429, n_1430, n_1431, n_1432, n_1433, n_1434, n_1435, n_1436, 
      n_1437, n_1438, n_1439, n_1440, n_1441, n_1442, n_1443, n_1444, n_1445, 
      n_1446, n_1447, n_1448, n_1449, n_1450, n_1451, n_1452, n_1453, n_1454, 
      n_1455, n_1456, n_1457, n_1458, n_1459, n_1460, n_1461, n_1462, n_1463, 
      n_1464, n_1465, n_1466, n_1467, n_1468, n_1469, n_1470, n_1471, n_1472, 
      n_1473, n_1474, n_1475, n_1476, n_1477, n_1478, n_1479, n_1480, n_1481, 
      n_1482, n_1483, n_1484, n_1485, n_1486, n_1487, n_1488, n_1489, n_1490, 
      n_1491, n_1492, n_1493, n_1494, n_1495, n_1496, n_1497, n_1498, n_1499, 
      n_1500, n_1501, n_1502, n_1503, n_1504, n_1505, n_1506, n_1507, n_1508, 
      n_1509, n_1510, n_1511, n_1512, n_1513, n_1514, n_1515, n_1516, n_1517, 
      n_1518, n_1519, n_1520, n_1521, n_1522, n_1523, n_1524, n_1525, n_1526, 
      n_1527, n_1528, n_1529, n_1530, n_1531, n_1532, n_1533, n_1534, n_1535, 
      n_1536, n_1537, n_1538, n_1539, n_1540, n_1541, n_1542, n_1543, n_1544, 
      n_1545, n_1546, n_1547, n_1548, n_1549, n_1550, n_1551, n_1552, n_1553, 
      n_1554, n_1555, n_1556, n_1557, n_1558, n_1559, n_1560, n_1561, n_1562, 
      n_1563, n_1564, n_1565, n_1566, n_1567, n_1568, n_1569, n_1570, n_1571, 
      n_1572, n_1573, n_1574, n_1575, n_1576, n_1577, n_1578, n_1579, n_1580, 
      n_1581, n_1582, n_1583, n_1584, n_1585, n_1586, n_1587, n_1588, n_1589, 
      n_1590, n_1591, n_1592, n_1593, n_1594, n_1595, n_1596, n_1597, n_1598, 
      n_1599, n_1600, n_1601, n_1602, n_1603, n_1604, n_1605, n_1606, n_1607, 
      n_1608, n_1609, n_1610, n_1611, n_1612, n_1613, n_1614, n_1615, n_1616, 
      n_1617, n_1618, n_1619, n_1620, n_1621, n_1622, n_1623, n_1624, n_1625, 
      n_1626, n_1627, n_1628, n_1629, n_1630, n_1631, n_1632, n_1633, n_1634, 
      n_1635, n_1636, n_1637, n_1638, n_1639, n_1640, n_1641, n_1642, n_1643, 
      n_1644, n_1645, n_1646, n_1647, n_1648, n_1649, n_1650, n_1651, n_1652, 
      n_1653, n_1654, n_1655, n_1656, n_1657, n_1658, n_1659, n_1660, n_1661, 
      n_1662, n_1663, n_1664, n_1665, n_1666, n_1667, n_1668, n_1669, n_1670, 
      n_1671, n_1672, n_1673, n_1674, n_1675, n_1676, n_1677, n_1678, n_1679, 
      n_1680, n_1681, n_1682, n_1683, n_1684, n_1685, n_1686, n_1687, n_1688, 
      n_1689, n_1690, n_1691, n_1692, n_1693, n_1694, n_1695, n_1696, n_1697, 
      n_1698, n_1699, n_1700, n_1701, n_1702, n_1703, n_1704, n_1705, n_1706, 
      n_1707, n_1708, n_1709, n_1710, n_1711, n_1712, n_1713, n_1714, n_1715, 
      n_1716, n_1717, n_1718, n_1719, n_1720, n_1721, n_1722, n_1723, n_1724, 
      n_1725, n_1726, n_1727, n_1728, n_1729, n_1730, n_1731, n_1732, n_1733, 
      n_1734, n_1735, n_1736, n_1737, n_1738, n_1739, n_1740, n_1741, n_1742, 
      n_1743, n_1744, n_1745, n_1746, n_1747, n_1748, n_1749, n_1750, n_1751, 
      n_1752, n_1753, n_1754, n_1755, n_1756, n_1757, n_1758, n_1759, n_1760, 
      n_1761, n_1762, n_1763, n_1764, n_1765, n_1766, n_1767, n_1768, n_1769, 
      n_1770, n_1771, n_1772, n_1773, n_1774, n_1775, n_1776, n_1777, n_1778, 
      n_1779, n_1780, n_1781, n_1782, n_1783, n_1784, n_1785, n_1786, n_1787, 
      n_1788, n_1789, n_1790, n_1791, n_1792, n_1793, n_1794, n_1795, n_1796, 
      n_1797, n_1798, n_1799, n_1800, n_1801, n_1802, n_1803, n_1804, n_1805, 
      n_1806, n_1807, n_1808, n_1809, n_1810, n_1811, n_1812, n_1813, n_1814, 
      n_1815, n_1816, n_1817, n_1818, n_1819, n_1820, n_1821, n_1822, n_1823, 
      n_1824, n_1825, n_1826, n_1827, n_1828, n_1829, n_1830, n_1831, n_1832, 
      n_1833, n_1834, n_1835, n_1836, n_1837, n_1838, n_1839, n_1840, n_1841, 
      n_1842, n_1843, n_1844, n_1845, n_1846, n_1847, n_1848, n_1849, n_1850, 
      n_1851, n_1852, n_1853, n_1854, n_1855, n_1856, n_1857, n_1858, n_1859, 
      n_1860, n_1861, n_1862, n_1863, n_1864, n_1865, n_1866, n_1867, n_1868, 
      n_1869, n_1870, n_1871, n_1872, n_1873, n_1874, n_1875, n_1876, n_1877, 
      n_1878, n_1879, n_1880, n_1881, n_1882, n_1883, n_1884, n_1885, n_1886, 
      n_1887, n_1888, n_1889, n_1890, n_1891, n_1892, n_1893, n_1894, n_1895, 
      n_1896, n_1897, n_1898, n_1899, n_1900, n_1901, n_1902, n_1903, n_1904, 
      n_1905, n_1906, n_1907, n_1908, n_1909, n_1910, n_1911, n_1912, n_1913, 
      n_1914, n_1915, n_1916, n_1917, n_1918, n_1919, n_1920, n_1921, n_1922, 
      n_1923, n_1924, n_1925, n_1926, n_1927, n_1928, n_1929, n_1930, n_1931, 
      n_1932, n_1933, n_1934, n_1935, n_1936, n_1937, n_1938, n_1939, n_1940, 
      n_1941, n_1942, n_1943, n_1944, n_1945, n_1946, n_1947, n_1948, n_1949, 
      n_1950, n_1951, n_1952, n_1953, n_1954, n_1955, n_1956, n_1957, n_1958, 
      n_1959, n_1960, n_1961, n_1962, n_1963, n_1964, n_1965, n_1966, n_1967, 
      n_1968, n_1969, n_1970, n_1971, n_1972, n_1973, n_1974, n_1975, n_1976, 
      n_1977, n_1978, n_1979, n_1980, n_1981, n_1982, n_1983, n_1984, n_1985, 
      n_1986, n_1987, n_1988, n_1989, n_1990, n_1991, n_1992, n_1993, n_1994, 
      n_1995, n_1996, n_1997, n_1998, n_1999, n_2000, n_2001, n_2002, n_2003, 
      n_2004, n_2005, n_2006, n_2007, n_2008, n_2009, n_2010, n_2011, n_2012, 
      n_2013, n_2014, n_2015, n_2016, n_2017, n_2018, n_2019, n_2020, n_2021, 
      n_2022, n_2023, n_2024, n_2025, n_2026, n_2027, n_2028, n_2029, n_2030, 
      n_2031, n_2032, n_2033, n_2034, n_2035, n_2036, n_2037, n_2038, n_2039, 
      n_2040, n_2041, n_2042, n_2043, n_2044, n_2045, n_2046, n_2047, n_2048, 
      n_2049, n_2050, n_2051, n_2052, n_2053, n_2054, n_2055, n_2056, n_2057, 
      n_2058, n_2059, n_2060, n_2061, n_2062, n_2063, n_2064, n_2065, n_2066, 
      n_2067, n_2068, n_2069, n_2070, n_2071, n_2072, n_2073, n_2074, n_2075, 
      n_2076, n_2077, n_2078, n_2079, n_2080, n_2081, n_2082, n_2083, n_2084, 
      n_2085, n_2086, n_2087, n_2088, n_2089, n_2090, n_2091, n_2092, n_2093, 
      n_2094, n_2095, n_2096, n_2097, n_2098, n_2099, n_2100, n_2101, n_2102, 
      n_2103, n_2104, n_2105, n_2106, n_2107, n_2108, n_2109, n_2110, n_2111, 
      n_2112, n_2113, n_2114, n_2115, n_2116, n_2117, n_2118, n_2119, n_2120, 
      n_2121, n_2122, n_2123, n_2124, n_2125, n_2126, n_2127, n_2128, n_2129, 
      n_2130, n_2131, n_2132, n_2133, n_2134, n_2135, n_2136, n_2137, n_2138, 
      n_2139, n_2140, n_2141, n_2142, n_2143, n_2144, n_2145, n_2146, n_2147, 
      n_2148, n_2149, n_2150, n_2151, n_2152, n_2153, n_2154, n_2155, n_2156, 
      n_2157, n_2158, n_2159, n_2160, n_2161, n_2162, n_2163, n_2164, n_2165, 
      n_2166, n_2167, n_2168, n_2169, n_2170, n_2171, n_2172, n_2173, n_2174, 
      n_2175, n_2176, n_2177, n_2178, n_2179, n_2180, n_2181, n_2182, n_2183, 
      n_2184, n_2185, n_2186, n_2187, n_2188, n_2189, n_2190, n_2191, n_2192, 
      n_2193, n_2194, n_2195, n_2196, n_2197, n_2198, n_2199, n_2200, n_2201, 
      n_2202, n_2203, n_2204, n_2205, n_2206, n_2207, n_2208, n_2209, n_2210, 
      n_2211 : std_logic;

begin
   
   n7 <= '0';
   n11 <= '0';
   n17 <= '0';
   REGISTERS_reg_0_31_inst : DFFR_X1 port map( D => n6317, CK => CLK, RN => 
                           n2974, Q => n3393, QN => n80);
   REGISTERS_reg_0_30_inst : DFFR_X1 port map( D => n6318, CK => CLK, RN => 
                           n2973, Q => n3395, QN => n81);
   REGISTERS_reg_0_29_inst : DFFR_X1 port map( D => n6319, CK => CLK, RN => 
                           n2971, Q => n3396, QN => n82);
   REGISTERS_reg_0_28_inst : DFFR_X1 port map( D => n6320, CK => CLK, RN => 
                           n2972, Q => n3397, QN => n83);
   REGISTERS_reg_0_27_inst : DFFR_X1 port map( D => n6321, CK => CLK, RN => 
                           n3264, Q => n3399, QN => n84);
   REGISTERS_reg_0_26_inst : DFFR_X1 port map( D => n6322, CK => CLK, RN => 
                           n3264, Q => n3401, QN => n85);
   REGISTERS_reg_0_25_inst : DFFR_X1 port map( D => n6323, CK => CLK, RN => 
                           n3264, Q => n3402, QN => n86);
   REGISTERS_reg_0_24_inst : DFFR_X1 port map( D => n6324, CK => CLK, RN => 
                           n3264, Q => n3404, QN => n87);
   REGISTERS_reg_0_23_inst : DFFR_X1 port map( D => n6325, CK => CLK, RN => 
                           n3264, Q => n3407, QN => n88);
   REGISTERS_reg_0_22_inst : DFFR_X1 port map( D => n6326, CK => CLK, RN => 
                           n3264, Q => n3408, QN => n89);
   REGISTERS_reg_0_21_inst : DFFR_X1 port map( D => n6327, CK => CLK, RN => 
                           n3264, Q => n3410, QN => n90);
   REGISTERS_reg_0_20_inst : DFFR_X1 port map( D => n6328, CK => CLK, RN => 
                           n3264, Q => n3411, QN => n91);
   REGISTERS_reg_0_19_inst : DFFR_X1 port map( D => n6329, CK => CLK, RN => 
                           n3264, Q => n3412, QN => n92);
   REGISTERS_reg_0_18_inst : DFFR_X1 port map( D => n6330, CK => CLK, RN => 
                           n3264, Q => n3414, QN => n93);
   REGISTERS_reg_0_17_inst : DFFR_X1 port map( D => n6331, CK => CLK, RN => 
                           n3264, Q => n9140, QN => n94);
   REGISTERS_reg_0_16_inst : DFFR_X1 port map( D => n6332, CK => CLK, RN => 
                           n3264, Q => n9141, QN => n95);
   REGISTERS_reg_0_15_inst : DFFR_X1 port map( D => n6333, CK => CLK, RN => 
                           n3262, Q => n9142, QN => n96);
   REGISTERS_reg_0_14_inst : DFFR_X1 port map( D => n6334, CK => CLK, RN => 
                           n3262, Q => n9143, QN => n97);
   REGISTERS_reg_0_13_inst : DFFR_X1 port map( D => n6335, CK => CLK, RN => 
                           n3262, Q => n9144, QN => n98);
   REGISTERS_reg_0_12_inst : DFFR_X1 port map( D => n6336, CK => CLK, RN => 
                           n3262, Q => n9145, QN => n99);
   REGISTERS_reg_0_11_inst : DFFR_X1 port map( D => n6337, CK => CLK, RN => 
                           n3262, Q => n9146, QN => n100);
   REGISTERS_reg_0_10_inst : DFFR_X1 port map( D => n6338, CK => CLK, RN => 
                           n3262, Q => n9147, QN => n101);
   REGISTERS_reg_0_9_inst : DFFR_X1 port map( D => n6339, CK => CLK, RN => 
                           n3262, Q => n9148, QN => n102);
   REGISTERS_reg_0_8_inst : DFFR_X1 port map( D => n6340, CK => CLK, RN => 
                           n3262, Q => n9149, QN => n103);
   REGISTERS_reg_0_7_inst : DFFR_X1 port map( D => n6341, CK => CLK, RN => 
                           n3262, Q => n9150, QN => n104);
   REGISTERS_reg_0_6_inst : DFFR_X1 port map( D => n6342, CK => CLK, RN => 
                           n3262, Q => n9151, QN => n105);
   REGISTERS_reg_0_5_inst : DFFR_X1 port map( D => n6343, CK => CLK, RN => 
                           n3262, Q => n9152, QN => n106);
   REGISTERS_reg_0_4_inst : DFFR_X1 port map( D => n6344, CK => CLK, RN => 
                           n3262, Q => n9153, QN => n107);
   REGISTERS_reg_0_3_inst : DFFR_X1 port map( D => n6345, CK => CLK, RN => 
                           n2977, Q => n9154, QN => n108);
   REGISTERS_reg_0_2_inst : DFFR_X1 port map( D => n6346, CK => CLK, RN => 
                           n2975, Q => n9155, QN => n109);
   REGISTERS_reg_0_1_inst : DFFR_X1 port map( D => n6347, CK => CLK, RN => 
                           n2976, Q => n9156, QN => n110);
   REGISTERS_reg_0_0_inst : DFFR_X1 port map( D => n6348, CK => CLK, RN => 
                           n3006, Q => n9157, QN => n111);
   REGISTERS_reg_1_31_inst : DFFR_X1 port map( D => n6349, CK => CLK, RN => 
                           n3007, Q => n9158, QN => n112);
   REGISTERS_reg_1_30_inst : DFFR_X1 port map( D => n6350, CK => CLK, RN => 
                           n2983, Q => n9159, QN => n113);
   REGISTERS_reg_1_29_inst : DFFR_X1 port map( D => n6351, CK => CLK, RN => 
                           n2981, Q => n9160, QN => n114);
   REGISTERS_reg_1_28_inst : DFFR_X1 port map( D => n6352, CK => CLK, RN => 
                           n2982, Q => n9161, QN => n115);
   REGISTERS_reg_1_27_inst : DFFR_X1 port map( D => n6353, CK => CLK, RN => 
                           n2984, Q => n9162, QN => n116);
   REGISTERS_reg_1_26_inst : DFFR_X1 port map( D => n6354, CK => CLK, RN => 
                           n2979, Q => n9163, QN => n117);
   REGISTERS_reg_1_25_inst : DFFR_X1 port map( D => n6355, CK => CLK, RN => 
                           n2980, Q => n9164, QN => n118);
   REGISTERS_reg_1_24_inst : DFFR_X1 port map( D => n6356, CK => CLK, RN => 
                           n2978, Q => n9165, QN => n119);
   REGISTERS_reg_1_23_inst : DFFR_X1 port map( D => n6357, CK => CLK, RN => 
                           n3018, Q => n9166, QN => n120);
   REGISTERS_reg_1_22_inst : DFFR_X1 port map( D => n6358, CK => CLK, RN => 
                           n3016, Q => n9167, QN => n121);
   REGISTERS_reg_1_21_inst : DFFR_X1 port map( D => n6359, CK => CLK, RN => 
                           n3014, Q => n9168, QN => n122);
   REGISTERS_reg_1_20_inst : DFFR_X1 port map( D => n6360, CK => CLK, RN => 
                           n3010, Q => n9169, QN => n123);
   REGISTERS_reg_1_19_inst : DFFR_X1 port map( D => n6361, CK => CLK, RN => 
                           n3017, Q => n9170, QN => n124);
   REGISTERS_reg_1_18_inst : DFFR_X1 port map( D => n6362, CK => CLK, RN => 
                           n3015, Q => n9171, QN => n125);
   REGISTERS_reg_1_17_inst : DFFR_X1 port map( D => n6363, CK => CLK, RN => 
                           n3011, Q => n9172, QN => n126);
   REGISTERS_reg_1_16_inst : DFFR_X1 port map( D => n6364, CK => CLK, RN => 
                           n3008, Q => n9173, QN => n127);
   REGISTERS_reg_1_15_inst : DFFR_X1 port map( D => n6365, CK => CLK, RN => 
                           n3019, Q => n9174, QN => n128);
   REGISTERS_reg_1_14_inst : DFFR_X1 port map( D => n6366, CK => CLK, RN => 
                           n3012, Q => n9175, QN => n129);
   REGISTERS_reg_1_13_inst : DFFR_X1 port map( D => n6367, CK => CLK, RN => 
                           n3013, Q => n9176, QN => n130);
   REGISTERS_reg_1_12_inst : DFFR_X1 port map( D => n6368, CK => CLK, RN => 
                           n3009, Q => n9177, QN => n131);
   REGISTERS_reg_1_11_inst : DFFR_X1 port map( D => n6369, CK => CLK, RN => 
                           n2990, Q => n9178, QN => n132);
   REGISTERS_reg_1_10_inst : DFFR_X1 port map( D => n6370, CK => CLK, RN => 
                           n2985, Q => n9179, QN => n133);
   REGISTERS_reg_1_9_inst : DFFR_X1 port map( D => n6371, CK => CLK, RN => 
                           n2986, Q => n9180, QN => n134);
   REGISTERS_reg_1_8_inst : DFFR_X1 port map( D => n6372, CK => CLK, RN => 
                           n3025, Q => n9181, QN => n135);
   REGISTERS_reg_1_7_inst : DFFR_X1 port map( D => n6373, CK => CLK, RN => 
                           n2989, Q => n9182, QN => n136);
   REGISTERS_reg_1_6_inst : DFFR_X1 port map( D => n6374, CK => CLK, RN => 
                           n2987, Q => n9183, QN => n137);
   REGISTERS_reg_1_5_inst : DFFR_X1 port map( D => n6375, CK => CLK, RN => 
                           n3023, Q => n9184, QN => n138);
   REGISTERS_reg_1_4_inst : DFFR_X1 port map( D => n6376, CK => CLK, RN => 
                           n3024, Q => n9185, QN => n139);
   REGISTERS_reg_1_3_inst : DFFR_X1 port map( D => n6377, CK => CLK, RN => 
                           n3022, Q => n9186, QN => n140);
   REGISTERS_reg_1_2_inst : DFFR_X1 port map( D => n6378, CK => CLK, RN => 
                           n3020, Q => n9187, QN => n141);
   REGISTERS_reg_1_1_inst : DFFR_X1 port map( D => n6379, CK => CLK, RN => 
                           n3021, Q => n9188, QN => n142);
   REGISTERS_reg_1_0_inst : DFFR_X1 port map( D => n6380, CK => CLK, RN => 
                           n2988, Q => n9189, QN => n143);
   REGISTERS_reg_2_31_inst : DFFR_X1 port map( D => n6381, CK => CLK, RN => 
                           n3261, Q => n9190, QN => n144);
   REGISTERS_reg_2_30_inst : DFFR_X1 port map( D => n6382, CK => CLK, RN => 
                           n3261, Q => n9191, QN => n145);
   REGISTERS_reg_2_29_inst : DFFR_X1 port map( D => n6383, CK => CLK, RN => 
                           n3261, Q => n9192, QN => n146);
   REGISTERS_reg_2_28_inst : DFFR_X1 port map( D => n6384, CK => CLK, RN => 
                           n3261, Q => n9193, QN => n147);
   REGISTERS_reg_2_27_inst : DFFR_X1 port map( D => n6385, CK => CLK, RN => 
                           n3261, Q => n9194, QN => n148);
   REGISTERS_reg_2_26_inst : DFFR_X1 port map( D => n6386, CK => CLK, RN => 
                           n3261, Q => n9195, QN => n149);
   REGISTERS_reg_2_25_inst : DFFR_X1 port map( D => n6387, CK => CLK, RN => 
                           n3261, Q => n9196, QN => n150);
   REGISTERS_reg_2_24_inst : DFFR_X1 port map( D => n6388, CK => CLK, RN => 
                           n3261, Q => n9197, QN => n151);
   REGISTERS_reg_2_23_inst : DFFR_X1 port map( D => n6389, CK => CLK, RN => 
                           n3261, Q => n9198, QN => n152);
   REGISTERS_reg_2_22_inst : DFFR_X1 port map( D => n6390, CK => CLK, RN => 
                           n3261, Q => n9199, QN => n153);
   REGISTERS_reg_2_21_inst : DFFR_X1 port map( D => n6391, CK => CLK, RN => 
                           n3261, Q => n9200, QN => n154);
   REGISTERS_reg_2_20_inst : DFFR_X1 port map( D => n6392, CK => CLK, RN => 
                           n3261, Q => n9201, QN => n155);
   REGISTERS_reg_2_19_inst : DFFR_X1 port map( D => n6393, CK => CLK, RN => 
                           n3260, Q => n9202, QN => n156);
   REGISTERS_reg_2_18_inst : DFFR_X1 port map( D => n6394, CK => CLK, RN => 
                           n3260, Q => n9203, QN => n157);
   REGISTERS_reg_2_17_inst : DFFR_X1 port map( D => n6395, CK => CLK, RN => 
                           n3260, Q => n9204, QN => n158);
   REGISTERS_reg_2_16_inst : DFFR_X1 port map( D => n6396, CK => CLK, RN => 
                           n3260, Q => n9205, QN => n159);
   REGISTERS_reg_2_15_inst : DFFR_X1 port map( D => n6397, CK => CLK, RN => 
                           n3260, Q => n9206, QN => n160);
   REGISTERS_reg_2_14_inst : DFFR_X1 port map( D => n6398, CK => CLK, RN => 
                           n3260, Q => n9207, QN => n161);
   REGISTERS_reg_2_13_inst : DFFR_X1 port map( D => n6399, CK => CLK, RN => 
                           n3260, Q => n9208, QN => n162);
   REGISTERS_reg_2_12_inst : DFFR_X1 port map( D => n6400, CK => CLK, RN => 
                           n3260, Q => n9209, QN => n163);
   REGISTERS_reg_2_11_inst : DFFR_X1 port map( D => n6401, CK => CLK, RN => 
                           n3260, Q => n9210, QN => n164);
   REGISTERS_reg_2_10_inst : DFFR_X1 port map( D => n6402, CK => CLK, RN => 
                           n3260, Q => n9211, QN => n165);
   REGISTERS_reg_2_9_inst : DFFR_X1 port map( D => n6403, CK => CLK, RN => 
                           n3260, Q => n9212, QN => n166);
   REGISTERS_reg_2_8_inst : DFFR_X1 port map( D => n6404, CK => CLK, RN => 
                           n3260, Q => n9213, QN => n167);
   REGISTERS_reg_2_7_inst : DFFR_X1 port map( D => n6405, CK => CLK, RN => 
                           n3258, Q => n9214, QN => n168);
   REGISTERS_reg_2_6_inst : DFFR_X1 port map( D => n6406, CK => CLK, RN => 
                           n3258, Q => n9215, QN => n169);
   REGISTERS_reg_2_5_inst : DFFR_X1 port map( D => n6407, CK => CLK, RN => 
                           n3258, Q => n9216, QN => n170);
   REGISTERS_reg_2_4_inst : DFFR_X1 port map( D => n6408, CK => CLK, RN => 
                           n3258, Q => n9217, QN => n171);
   REGISTERS_reg_2_3_inst : DFFR_X1 port map( D => n6409, CK => CLK, RN => 
                           n3258, Q => n9218, QN => n172);
   REGISTERS_reg_2_2_inst : DFFR_X1 port map( D => n6410, CK => CLK, RN => 
                           n3258, Q => n9219, QN => n173);
   REGISTERS_reg_2_1_inst : DFFR_X1 port map( D => n6411, CK => CLK, RN => 
                           n3258, Q => n9220, QN => n174);
   REGISTERS_reg_2_0_inst : DFFR_X1 port map( D => n6412, CK => CLK, RN => 
                           n3258, Q => n9221, QN => n175);
   REGISTERS_reg_3_31_inst : DFFR_X1 port map( D => n6413, CK => CLK, RN => 
                           n3258, Q => n9222, QN => n176);
   REGISTERS_reg_3_30_inst : DFFR_X1 port map( D => n6414, CK => CLK, RN => 
                           n3258, Q => n9223, QN => n177);
   REGISTERS_reg_3_29_inst : DFFR_X1 port map( D => n6415, CK => CLK, RN => 
                           n3258, Q => n9224, QN => n178);
   REGISTERS_reg_3_28_inst : DFFR_X1 port map( D => n6416, CK => CLK, RN => 
                           n3258, Q => n9225, QN => n179);
   REGISTERS_reg_3_27_inst : DFFR_X1 port map( D => n6417, CK => CLK, RN => 
                           n3257, Q => n9226, QN => n180);
   REGISTERS_reg_3_26_inst : DFFR_X1 port map( D => n6418, CK => CLK, RN => 
                           n3257, Q => n9227, QN => n181);
   REGISTERS_reg_3_25_inst : DFFR_X1 port map( D => n6419, CK => CLK, RN => 
                           n3257, Q => n9228, QN => n182);
   REGISTERS_reg_3_24_inst : DFFR_X1 port map( D => n6420, CK => CLK, RN => 
                           n3257, Q => n9229, QN => n183);
   REGISTERS_reg_3_23_inst : DFFR_X1 port map( D => n6421, CK => CLK, RN => 
                           n3257, Q => n9230, QN => n184);
   REGISTERS_reg_3_22_inst : DFFR_X1 port map( D => n6422, CK => CLK, RN => 
                           n3257, Q => n9231, QN => n185);
   REGISTERS_reg_3_21_inst : DFFR_X1 port map( D => n6423, CK => CLK, RN => 
                           n3257, Q => n9232, QN => n186);
   REGISTERS_reg_3_20_inst : DFFR_X1 port map( D => n6424, CK => CLK, RN => 
                           n3257, Q => n9233, QN => n187);
   REGISTERS_reg_3_19_inst : DFFR_X1 port map( D => n6425, CK => CLK, RN => 
                           n3257, Q => n9234, QN => n188);
   REGISTERS_reg_3_18_inst : DFFR_X1 port map( D => n6426, CK => CLK, RN => 
                           n3257, Q => n9235, QN => n189);
   REGISTERS_reg_3_17_inst : DFFR_X1 port map( D => n6427, CK => CLK, RN => 
                           n3257, Q => n9236, QN => n190);
   REGISTERS_reg_3_16_inst : DFFR_X1 port map( D => n6428, CK => CLK, RN => 
                           n3257, Q => n9237, QN => n191);
   REGISTERS_reg_3_15_inst : DFFR_X1 port map( D => n6429, CK => CLK, RN => 
                           n3256, Q => n9238, QN => n192);
   REGISTERS_reg_3_14_inst : DFFR_X1 port map( D => n6430, CK => CLK, RN => 
                           n3256, Q => n9239, QN => n193);
   REGISTERS_reg_3_13_inst : DFFR_X1 port map( D => n6431, CK => CLK, RN => 
                           n3256, Q => n9240, QN => n194);
   REGISTERS_reg_3_12_inst : DFFR_X1 port map( D => n6432, CK => CLK, RN => 
                           n3256, Q => n9241, QN => n195);
   REGISTERS_reg_3_11_inst : DFFR_X1 port map( D => n6433, CK => CLK, RN => 
                           n3256, Q => n9242, QN => n196);
   REGISTERS_reg_3_10_inst : DFFR_X1 port map( D => n6434, CK => CLK, RN => 
                           n3256, Q => n9243, QN => n197);
   REGISTERS_reg_3_9_inst : DFFR_X1 port map( D => n6435, CK => CLK, RN => 
                           n3256, Q => n9244, QN => n198);
   REGISTERS_reg_3_8_inst : DFFR_X1 port map( D => n6436, CK => CLK, RN => 
                           n3256, Q => n9245, QN => n199);
   REGISTERS_reg_3_7_inst : DFFR_X1 port map( D => n6437, CK => CLK, RN => 
                           n3256, Q => n9246, QN => n200);
   REGISTERS_reg_3_6_inst : DFFR_X1 port map( D => n6438, CK => CLK, RN => 
                           n3256, Q => n9247, QN => n201);
   REGISTERS_reg_3_5_inst : DFFR_X1 port map( D => n6439, CK => CLK, RN => 
                           n3256, Q => n9248, QN => n202);
   REGISTERS_reg_3_4_inst : DFFR_X1 port map( D => n6440, CK => CLK, RN => 
                           n3256, Q => n9249, QN => n203);
   REGISTERS_reg_3_3_inst : DFFR_X1 port map( D => n6441, CK => CLK, RN => 
                           n3254, Q => n9250, QN => n204);
   REGISTERS_reg_3_2_inst : DFFR_X1 port map( D => n6442, CK => CLK, RN => 
                           n3254, Q => n9251, QN => n205);
   REGISTERS_reg_3_1_inst : DFFR_X1 port map( D => n6443, CK => CLK, RN => 
                           n3254, Q => n9252, QN => n206);
   REGISTERS_reg_3_0_inst : DFFR_X1 port map( D => n6444, CK => CLK, RN => 
                           n3254, Q => n9253, QN => n207);
   REGISTERS_reg_4_31_inst : DFFR_X1 port map( D => n6445, CK => CLK, RN => 
                           n3254, Q => n9254, QN => n208);
   REGISTERS_reg_4_30_inst : DFFR_X1 port map( D => n6446, CK => CLK, RN => 
                           n3254, Q => n9255, QN => n209);
   REGISTERS_reg_4_29_inst : DFFR_X1 port map( D => n6447, CK => CLK, RN => 
                           n3254, Q => n9256, QN => n210);
   REGISTERS_reg_4_28_inst : DFFR_X1 port map( D => n6448, CK => CLK, RN => 
                           n3254, Q => n9257, QN => n211);
   REGISTERS_reg_4_27_inst : DFFR_X1 port map( D => n6449, CK => CLK, RN => 
                           n3254, Q => n9258, QN => n212);
   REGISTERS_reg_4_26_inst : DFFR_X1 port map( D => n6450, CK => CLK, RN => 
                           n3254, Q => n9259, QN => n213);
   REGISTERS_reg_4_25_inst : DFFR_X1 port map( D => n6451, CK => CLK, RN => 
                           n3254, Q => n9260, QN => n214);
   REGISTERS_reg_4_24_inst : DFFR_X1 port map( D => n6452, CK => CLK, RN => 
                           n3254, Q => n9261, QN => n215);
   REGISTERS_reg_4_23_inst : DFFR_X1 port map( D => n6453, CK => CLK, RN => 
                           n3253, Q => n9262, QN => n216);
   REGISTERS_reg_4_22_inst : DFFR_X1 port map( D => n6454, CK => CLK, RN => 
                           n3253, Q => n9263, QN => n217);
   REGISTERS_reg_4_21_inst : DFFR_X1 port map( D => n6455, CK => CLK, RN => 
                           n3253, Q => n9264, QN => n218);
   REGISTERS_reg_4_20_inst : DFFR_X1 port map( D => n6456, CK => CLK, RN => 
                           n3253, Q => n9265, QN => n219);
   REGISTERS_reg_4_19_inst : DFFR_X1 port map( D => n6457, CK => CLK, RN => 
                           n3253, Q => n9266, QN => n220);
   REGISTERS_reg_4_18_inst : DFFR_X1 port map( D => n6458, CK => CLK, RN => 
                           n3253, Q => n9267, QN => n221);
   REGISTERS_reg_4_17_inst : DFFR_X1 port map( D => n6459, CK => CLK, RN => 
                           n3253, Q => n9268, QN => n222);
   REGISTERS_reg_4_16_inst : DFFR_X1 port map( D => n6460, CK => CLK, RN => 
                           n3253, Q => n9269, QN => n223);
   REGISTERS_reg_4_15_inst : DFFR_X1 port map( D => n6461, CK => CLK, RN => 
                           n3253, Q => n9270, QN => n224);
   REGISTERS_reg_4_14_inst : DFFR_X1 port map( D => n6462, CK => CLK, RN => 
                           n3253, Q => n9271, QN => n225);
   REGISTERS_reg_4_13_inst : DFFR_X1 port map( D => n6463, CK => CLK, RN => 
                           n3253, Q => n9272, QN => n226);
   REGISTERS_reg_4_12_inst : DFFR_X1 port map( D => n6464, CK => CLK, RN => 
                           n3253, Q => n9273, QN => n227);
   REGISTERS_reg_4_11_inst : DFFR_X1 port map( D => n6465, CK => CLK, RN => 
                           n3252, Q => n9274, QN => n228);
   REGISTERS_reg_4_10_inst : DFFR_X1 port map( D => n6466, CK => CLK, RN => 
                           n3252, Q => n9275, QN => n229);
   REGISTERS_reg_4_9_inst : DFFR_X1 port map( D => n6467, CK => CLK, RN => 
                           n3252, Q => n9276, QN => n230);
   REGISTERS_reg_4_8_inst : DFFR_X1 port map( D => n6468, CK => CLK, RN => 
                           n3252, Q => n9277, QN => n231);
   REGISTERS_reg_4_7_inst : DFFR_X1 port map( D => n6469, CK => CLK, RN => 
                           n3252, Q => n9278, QN => n232);
   REGISTERS_reg_4_6_inst : DFFR_X1 port map( D => n6470, CK => CLK, RN => 
                           n3252, Q => n9279, QN => n233);
   REGISTERS_reg_4_5_inst : DFFR_X1 port map( D => n6471, CK => CLK, RN => 
                           n3252, Q => n9280, QN => n234);
   REGISTERS_reg_4_4_inst : DFFR_X1 port map( D => n6472, CK => CLK, RN => 
                           n3252, Q => n9281, QN => n235);
   REGISTERS_reg_4_3_inst : DFFR_X1 port map( D => n6473, CK => CLK, RN => 
                           n3252, Q => n9282, QN => n236);
   REGISTERS_reg_4_2_inst : DFFR_X1 port map( D => n6474, CK => CLK, RN => 
                           n3252, Q => n9283, QN => n237);
   REGISTERS_reg_4_1_inst : DFFR_X1 port map( D => n6475, CK => CLK, RN => 
                           n3252, Q => n9284, QN => n238);
   REGISTERS_reg_4_0_inst : DFFR_X1 port map( D => n6476, CK => CLK, RN => 
                           n3252, Q => n9285, QN => n239);
   REGISTERS_reg_5_31_inst : DFFR_X1 port map( D => n6477, CK => CLK, RN => 
                           n3250, Q => n9286, QN => n240);
   REGISTERS_reg_5_30_inst : DFFR_X1 port map( D => n6478, CK => CLK, RN => 
                           n3250, Q => n9287, QN => n241);
   REGISTERS_reg_5_29_inst : DFFR_X1 port map( D => n6479, CK => CLK, RN => 
                           n3250, Q => n9288, QN => n242);
   REGISTERS_reg_5_28_inst : DFFR_X1 port map( D => n6480, CK => CLK, RN => 
                           n3250, Q => n9289, QN => n243);
   REGISTERS_reg_5_27_inst : DFFR_X1 port map( D => n6481, CK => CLK, RN => 
                           n3250, Q => n9290, QN => n244);
   REGISTERS_reg_5_26_inst : DFFR_X1 port map( D => n6482, CK => CLK, RN => 
                           n3250, Q => n9291, QN => n245);
   REGISTERS_reg_5_25_inst : DFFR_X1 port map( D => n6483, CK => CLK, RN => 
                           n3250, Q => n9292, QN => n246);
   REGISTERS_reg_5_24_inst : DFFR_X1 port map( D => n6484, CK => CLK, RN => 
                           n3250, Q => n9293, QN => n247);
   REGISTERS_reg_5_23_inst : DFFR_X1 port map( D => n6485, CK => CLK, RN => 
                           n3250, Q => n9294, QN => n248);
   REGISTERS_reg_5_22_inst : DFFR_X1 port map( D => n6486, CK => CLK, RN => 
                           n3250, Q => n9295, QN => n249);
   REGISTERS_reg_5_21_inst : DFFR_X1 port map( D => n6487, CK => CLK, RN => 
                           n3250, Q => n9296, QN => n250);
   REGISTERS_reg_5_20_inst : DFFR_X1 port map( D => n6488, CK => CLK, RN => 
                           n3250, Q => n9297, QN => n251);
   REGISTERS_reg_5_19_inst : DFFR_X1 port map( D => n6489, CK => CLK, RN => 
                           n3249, Q => n9298, QN => n252);
   REGISTERS_reg_5_18_inst : DFFR_X1 port map( D => n6490, CK => CLK, RN => 
                           n3249, Q => n9299, QN => n253);
   REGISTERS_reg_5_17_inst : DFFR_X1 port map( D => n6491, CK => CLK, RN => 
                           n3249, Q => n9300, QN => n254);
   REGISTERS_reg_5_16_inst : DFFR_X1 port map( D => n6492, CK => CLK, RN => 
                           n3249, Q => n9301, QN => n255);
   REGISTERS_reg_5_15_inst : DFFR_X1 port map( D => n6493, CK => CLK, RN => 
                           n3249, Q => n9302, QN => n256);
   REGISTERS_reg_5_14_inst : DFFR_X1 port map( D => n6494, CK => CLK, RN => 
                           n3249, Q => n9303, QN => n257);
   REGISTERS_reg_5_13_inst : DFFR_X1 port map( D => n6495, CK => CLK, RN => 
                           n3249, Q => n9304, QN => n258);
   REGISTERS_reg_5_12_inst : DFFR_X1 port map( D => n6496, CK => CLK, RN => 
                           n3249, Q => n9305, QN => n259);
   REGISTERS_reg_5_11_inst : DFFR_X1 port map( D => n6497, CK => CLK, RN => 
                           n3249, Q => n9306, QN => n260);
   REGISTERS_reg_5_10_inst : DFFR_X1 port map( D => n6498, CK => CLK, RN => 
                           n3249, Q => n9307, QN => n261);
   REGISTERS_reg_5_9_inst : DFFR_X1 port map( D => n6499, CK => CLK, RN => 
                           n3249, Q => n9308, QN => n262);
   REGISTERS_reg_5_8_inst : DFFR_X1 port map( D => n6500, CK => CLK, RN => 
                           n3249, Q => n9309, QN => n263);
   REGISTERS_reg_5_7_inst : DFFR_X1 port map( D => n6501, CK => CLK, RN => 
                           n3248, Q => n9310, QN => n264);
   REGISTERS_reg_5_6_inst : DFFR_X1 port map( D => n6502, CK => CLK, RN => 
                           n3248, Q => n9311, QN => n265);
   REGISTERS_reg_5_5_inst : DFFR_X1 port map( D => n6503, CK => CLK, RN => 
                           n3248, Q => n9312, QN => n266);
   REGISTERS_reg_5_4_inst : DFFR_X1 port map( D => n6504, CK => CLK, RN => 
                           n3248, Q => n9313, QN => n267);
   REGISTERS_reg_5_3_inst : DFFR_X1 port map( D => n6505, CK => CLK, RN => 
                           n3248, Q => n9314, QN => n268);
   REGISTERS_reg_5_2_inst : DFFR_X1 port map( D => n6506, CK => CLK, RN => 
                           n3248, Q => n9315, QN => n269);
   REGISTERS_reg_5_1_inst : DFFR_X1 port map( D => n6507, CK => CLK, RN => 
                           n3248, Q => n9316, QN => n270);
   REGISTERS_reg_5_0_inst : DFFR_X1 port map( D => n6508, CK => CLK, RN => 
                           n3248, Q => n9317, QN => n271);
   REGISTERS_reg_6_31_inst : DFFR_X1 port map( D => n6509, CK => CLK, RN => 
                           n3248, Q => n9318, QN => n272);
   REGISTERS_reg_6_30_inst : DFFR_X1 port map( D => n6510, CK => CLK, RN => 
                           n3248, Q => n9319, QN => n273);
   REGISTERS_reg_6_29_inst : DFFR_X1 port map( D => n6511, CK => CLK, RN => 
                           n3248, Q => n9320, QN => n274);
   REGISTERS_reg_6_28_inst : DFFR_X1 port map( D => n6512, CK => CLK, RN => 
                           n3248, Q => n9321, QN => n275);
   REGISTERS_reg_6_27_inst : DFFR_X1 port map( D => n6513, CK => CLK, RN => 
                           n3246, Q => n9322, QN => n276);
   REGISTERS_reg_6_26_inst : DFFR_X1 port map( D => n6514, CK => CLK, RN => 
                           n3246, Q => n9323, QN => n277);
   REGISTERS_reg_6_25_inst : DFFR_X1 port map( D => n6515, CK => CLK, RN => 
                           n3246, Q => n9324, QN => n278);
   REGISTERS_reg_6_24_inst : DFFR_X1 port map( D => n6516, CK => CLK, RN => 
                           n3246, Q => n9325, QN => n279);
   REGISTERS_reg_6_23_inst : DFFR_X1 port map( D => n6517, CK => CLK, RN => 
                           n3246, Q => n9326, QN => n280);
   REGISTERS_reg_6_22_inst : DFFR_X1 port map( D => n6518, CK => CLK, RN => 
                           n3246, Q => n9327, QN => n281);
   REGISTERS_reg_6_21_inst : DFFR_X1 port map( D => n6519, CK => CLK, RN => 
                           n3246, Q => n9328, QN => n282);
   REGISTERS_reg_6_20_inst : DFFR_X1 port map( D => n6520, CK => CLK, RN => 
                           n3246, Q => n9329, QN => n283);
   REGISTERS_reg_6_19_inst : DFFR_X1 port map( D => n6521, CK => CLK, RN => 
                           n3246, Q => n9330, QN => n284);
   REGISTERS_reg_6_18_inst : DFFR_X1 port map( D => n6522, CK => CLK, RN => 
                           n3246, Q => n9331, QN => n285);
   REGISTERS_reg_6_17_inst : DFFR_X1 port map( D => n6523, CK => CLK, RN => 
                           n3246, Q => n9332, QN => n286);
   REGISTERS_reg_6_16_inst : DFFR_X1 port map( D => n6524, CK => CLK, RN => 
                           n3246, Q => n9333, QN => n287);
   REGISTERS_reg_6_15_inst : DFFR_X1 port map( D => n6525, CK => CLK, RN => 
                           n3245, Q => n9334, QN => n288);
   REGISTERS_reg_6_14_inst : DFFR_X1 port map( D => n6526, CK => CLK, RN => 
                           n3245, Q => n9335, QN => n289);
   REGISTERS_reg_6_13_inst : DFFR_X1 port map( D => n6527, CK => CLK, RN => 
                           n3245, Q => n9336, QN => n290);
   REGISTERS_reg_6_12_inst : DFFR_X1 port map( D => n6528, CK => CLK, RN => 
                           n3245, Q => n9337, QN => n291);
   REGISTERS_reg_6_11_inst : DFFR_X1 port map( D => n6529, CK => CLK, RN => 
                           n3245, Q => n9338, QN => n292);
   REGISTERS_reg_6_10_inst : DFFR_X1 port map( D => n6530, CK => CLK, RN => 
                           n3245, Q => n9339, QN => n293);
   REGISTERS_reg_6_9_inst : DFFR_X1 port map( D => n6531, CK => CLK, RN => 
                           n3245, Q => n9340, QN => n294);
   REGISTERS_reg_6_8_inst : DFFR_X1 port map( D => n6532, CK => CLK, RN => 
                           n3245, Q => n9341, QN => n295);
   REGISTERS_reg_6_7_inst : DFFR_X1 port map( D => n6533, CK => CLK, RN => 
                           n3245, Q => n9342, QN => n296);
   REGISTERS_reg_6_6_inst : DFFR_X1 port map( D => n6534, CK => CLK, RN => 
                           n3245, Q => n9343, QN => n297);
   REGISTERS_reg_6_5_inst : DFFR_X1 port map( D => n6535, CK => CLK, RN => 
                           n3245, Q => n9344, QN => n298);
   REGISTERS_reg_6_4_inst : DFFR_X1 port map( D => n6536, CK => CLK, RN => 
                           n3245, Q => n9345, QN => n299);
   REGISTERS_reg_6_3_inst : DFFR_X1 port map( D => n6537, CK => CLK, RN => 
                           n3243, Q => n9346, QN => n300);
   REGISTERS_reg_6_2_inst : DFFR_X1 port map( D => n6538, CK => CLK, RN => 
                           n3243, Q => n9347, QN => n301);
   REGISTERS_reg_6_1_inst : DFFR_X1 port map( D => n6539, CK => CLK, RN => 
                           n3243, Q => n9348, QN => n302);
   REGISTERS_reg_6_0_inst : DFFR_X1 port map( D => n6540, CK => CLK, RN => 
                           n3243, Q => n9349, QN => n303);
   REGISTERS_reg_7_31_inst : DFFR_X1 port map( D => n6541, CK => CLK, RN => 
                           n3243, Q => n9350, QN => n304);
   REGISTERS_reg_7_30_inst : DFFR_X1 port map( D => n6542, CK => CLK, RN => 
                           n3243, Q => n9351, QN => n305);
   REGISTERS_reg_7_29_inst : DFFR_X1 port map( D => n6543, CK => CLK, RN => 
                           n3243, Q => n9352, QN => n306);
   REGISTERS_reg_7_28_inst : DFFR_X1 port map( D => n6544, CK => CLK, RN => 
                           n3243, Q => n9353, QN => n307);
   REGISTERS_reg_7_27_inst : DFFR_X1 port map( D => n6545, CK => CLK, RN => 
                           n3243, Q => n9354, QN => n308);
   REGISTERS_reg_7_26_inst : DFFR_X1 port map( D => n6546, CK => CLK, RN => 
                           n3243, Q => n9355, QN => n309);
   REGISTERS_reg_7_25_inst : DFFR_X1 port map( D => n6547, CK => CLK, RN => 
                           n3243, Q => n9356, QN => n310);
   REGISTERS_reg_7_24_inst : DFFR_X1 port map( D => n6548, CK => CLK, RN => 
                           n3243, Q => n9357, QN => n311);
   REGISTERS_reg_7_23_inst : DFFR_X1 port map( D => n6549, CK => CLK, RN => 
                           n3241, Q => n9358, QN => n312);
   REGISTERS_reg_7_22_inst : DFFR_X1 port map( D => n6550, CK => CLK, RN => 
                           n3241, Q => n9359, QN => n313);
   REGISTERS_reg_7_21_inst : DFFR_X1 port map( D => n6551, CK => CLK, RN => 
                           n3241, Q => n9360, QN => n314);
   REGISTERS_reg_7_20_inst : DFFR_X1 port map( D => n6552, CK => CLK, RN => 
                           n3241, Q => n9361, QN => n315);
   REGISTERS_reg_7_19_inst : DFFR_X1 port map( D => n6553, CK => CLK, RN => 
                           n3241, Q => n9362, QN => n316);
   REGISTERS_reg_7_18_inst : DFFR_X1 port map( D => n6554, CK => CLK, RN => 
                           n3241, Q => n9363, QN => n317);
   REGISTERS_reg_7_17_inst : DFFR_X1 port map( D => n6555, CK => CLK, RN => 
                           n3241, Q => n9364, QN => n318);
   REGISTERS_reg_7_16_inst : DFFR_X1 port map( D => n6556, CK => CLK, RN => 
                           n3241, Q => n9365, QN => n319);
   REGISTERS_reg_7_15_inst : DFFR_X1 port map( D => n6557, CK => CLK, RN => 
                           n3241, Q => n9366, QN => n320);
   REGISTERS_reg_7_14_inst : DFFR_X1 port map( D => n6558, CK => CLK, RN => 
                           n3241, Q => n9367, QN => n321);
   REGISTERS_reg_7_13_inst : DFFR_X1 port map( D => n6559, CK => CLK, RN => 
                           n3241, Q => n9368, QN => n322);
   REGISTERS_reg_7_12_inst : DFFR_X1 port map( D => n6560, CK => CLK, RN => 
                           n3241, Q => n9369, QN => n323);
   REGISTERS_reg_7_11_inst : DFFR_X1 port map( D => n6561, CK => CLK, RN => 
                           n3240, Q => n9370, QN => n324);
   REGISTERS_reg_7_10_inst : DFFR_X1 port map( D => n6562, CK => CLK, RN => 
                           n3240, Q => n9371, QN => n325);
   REGISTERS_reg_7_9_inst : DFFR_X1 port map( D => n6563, CK => CLK, RN => 
                           n3240, Q => n9372, QN => n326);
   REGISTERS_reg_7_8_inst : DFFR_X1 port map( D => n6564, CK => CLK, RN => 
                           n3240, Q => n9373, QN => n327);
   REGISTERS_reg_7_7_inst : DFFR_X1 port map( D => n6565, CK => CLK, RN => 
                           n3240, Q => n9374, QN => n328);
   REGISTERS_reg_7_6_inst : DFFR_X1 port map( D => n6566, CK => CLK, RN => 
                           n3240, Q => n9375, QN => n329);
   REGISTERS_reg_7_5_inst : DFFR_X1 port map( D => n6567, CK => CLK, RN => 
                           n3240, Q => n9376, QN => n330);
   REGISTERS_reg_7_4_inst : DFFR_X1 port map( D => n6568, CK => CLK, RN => 
                           n3240, Q => n9377, QN => n331);
   REGISTERS_reg_7_3_inst : DFFR_X1 port map( D => n6569, CK => CLK, RN => 
                           n3240, Q => n9378, QN => n332);
   REGISTERS_reg_7_2_inst : DFFR_X1 port map( D => n6570, CK => CLK, RN => 
                           n3240, Q => n9379, QN => n333);
   REGISTERS_reg_7_1_inst : DFFR_X1 port map( D => n6571, CK => CLK, RN => 
                           n3240, Q => n9380, QN => n334);
   REGISTERS_reg_7_0_inst : DFFR_X1 port map( D => n6572, CK => CLK, RN => 
                           n3240, Q => n9381, QN => n335);
   REGISTERS_reg_8_31_inst : DFFR_X1 port map( D => n6573, CK => CLK, RN => 
                           n3239, Q => n9382, QN => n336);
   REGISTERS_reg_8_30_inst : DFFR_X1 port map( D => n6574, CK => CLK, RN => 
                           n3239, Q => n9383, QN => n337);
   REGISTERS_reg_8_29_inst : DFFR_X1 port map( D => n6575, CK => CLK, RN => 
                           n3239, Q => n9384, QN => n338);
   REGISTERS_reg_8_28_inst : DFFR_X1 port map( D => n6576, CK => CLK, RN => 
                           n3239, Q => n9385, QN => n339);
   REGISTERS_reg_8_27_inst : DFFR_X1 port map( D => n6577, CK => CLK, RN => 
                           n3239, Q => n9386, QN => n340);
   REGISTERS_reg_8_26_inst : DFFR_X1 port map( D => n6578, CK => CLK, RN => 
                           n3239, Q => n9387, QN => n341);
   REGISTERS_reg_8_25_inst : DFFR_X1 port map( D => n6579, CK => CLK, RN => 
                           n3239, Q => n9388, QN => n342);
   REGISTERS_reg_8_24_inst : DFFR_X1 port map( D => n6580, CK => CLK, RN => 
                           n3239, Q => n9389, QN => n343);
   REGISTERS_reg_8_23_inst : DFFR_X1 port map( D => n6581, CK => CLK, RN => 
                           n3239, Q => n9390, QN => n344);
   REGISTERS_reg_8_22_inst : DFFR_X1 port map( D => n6582, CK => CLK, RN => 
                           n3239, Q => n9391, QN => n345);
   REGISTERS_reg_8_21_inst : DFFR_X1 port map( D => n6583, CK => CLK, RN => 
                           n3239, Q => n9392, QN => n346);
   REGISTERS_reg_8_20_inst : DFFR_X1 port map( D => n6584, CK => CLK, RN => 
                           n3239, Q => n9393, QN => n347);
   REGISTERS_reg_8_19_inst : DFFR_X1 port map( D => n6585, CK => CLK, RN => 
                           n3237, Q => n9394, QN => n348);
   REGISTERS_reg_8_18_inst : DFFR_X1 port map( D => n6586, CK => CLK, RN => 
                           n3237, Q => n9395, QN => n349);
   REGISTERS_reg_8_17_inst : DFFR_X1 port map( D => n6587, CK => CLK, RN => 
                           n3237, Q => n9396, QN => n350);
   REGISTERS_reg_8_16_inst : DFFR_X1 port map( D => n6588, CK => CLK, RN => 
                           n3237, Q => n9397, QN => n351);
   REGISTERS_reg_8_15_inst : DFFR_X1 port map( D => n6589, CK => CLK, RN => 
                           n3237, Q => n9398, QN => n352);
   REGISTERS_reg_8_14_inst : DFFR_X1 port map( D => n6590, CK => CLK, RN => 
                           n3237, Q => n9399, QN => n353);
   REGISTERS_reg_8_13_inst : DFFR_X1 port map( D => n6591, CK => CLK, RN => 
                           n3237, Q => n9400, QN => n354);
   REGISTERS_reg_8_12_inst : DFFR_X1 port map( D => n6592, CK => CLK, RN => 
                           n3237, Q => n9401, QN => n355);
   REGISTERS_reg_8_11_inst : DFFR_X1 port map( D => n6593, CK => CLK, RN => 
                           n3237, Q => n9402, QN => n356);
   REGISTERS_reg_8_10_inst : DFFR_X1 port map( D => n6594, CK => CLK, RN => 
                           n3237, Q => n9403, QN => n357);
   REGISTERS_reg_8_9_inst : DFFR_X1 port map( D => n6595, CK => CLK, RN => 
                           n3237, Q => n9404, QN => n358);
   REGISTERS_reg_8_8_inst : DFFR_X1 port map( D => n6596, CK => CLK, RN => 
                           n3237, Q => n9405, QN => n359);
   REGISTERS_reg_8_7_inst : DFFR_X1 port map( D => n6597, CK => CLK, RN => 
                           n3236, Q => n9406, QN => n360);
   REGISTERS_reg_8_6_inst : DFFR_X1 port map( D => n6598, CK => CLK, RN => 
                           n3236, Q => n9407, QN => n361);
   REGISTERS_reg_8_5_inst : DFFR_X1 port map( D => n6599, CK => CLK, RN => 
                           n3236, Q => n9408, QN => n362);
   REGISTERS_reg_8_4_inst : DFFR_X1 port map( D => n6600, CK => CLK, RN => 
                           n3236, Q => n9409, QN => n363);
   REGISTERS_reg_8_3_inst : DFFR_X1 port map( D => n6601, CK => CLK, RN => 
                           n3236, Q => n9410, QN => n364);
   REGISTERS_reg_8_2_inst : DFFR_X1 port map( D => n6602, CK => CLK, RN => 
                           n3236, Q => n9411, QN => n365);
   REGISTERS_reg_8_1_inst : DFFR_X1 port map( D => n6603, CK => CLK, RN => 
                           n3236, Q => n9412, QN => n366);
   REGISTERS_reg_8_0_inst : DFFR_X1 port map( D => n6604, CK => CLK, RN => 
                           n3236, Q => n9413, QN => n367);
   REGISTERS_reg_9_31_inst : DFFR_X1 port map( D => n6605, CK => CLK, RN => 
                           n3236, Q => n9414, QN => n368);
   REGISTERS_reg_9_30_inst : DFFR_X1 port map( D => n6606, CK => CLK, RN => 
                           n3236, Q => n9415, QN => n369);
   REGISTERS_reg_9_29_inst : DFFR_X1 port map( D => n6607, CK => CLK, RN => 
                           n3236, Q => n9416, QN => n370);
   REGISTERS_reg_9_28_inst : DFFR_X1 port map( D => n6608, CK => CLK, RN => 
                           n3236, Q => n9417, QN => n371);
   REGISTERS_reg_9_27_inst : DFFR_X1 port map( D => n6609, CK => CLK, RN => 
                           n3235, Q => n9418, QN => n372);
   REGISTERS_reg_9_26_inst : DFFR_X1 port map( D => n6610, CK => CLK, RN => 
                           n3235, Q => n9419, QN => n373);
   REGISTERS_reg_9_25_inst : DFFR_X1 port map( D => n6611, CK => CLK, RN => 
                           n3235, Q => n9420, QN => n374);
   REGISTERS_reg_9_24_inst : DFFR_X1 port map( D => n6612, CK => CLK, RN => 
                           n3235, Q => n9421, QN => n375);
   REGISTERS_reg_9_23_inst : DFFR_X1 port map( D => n6613, CK => CLK, RN => 
                           n3235, Q => n9422, QN => n376);
   REGISTERS_reg_9_22_inst : DFFR_X1 port map( D => n6614, CK => CLK, RN => 
                           n3235, Q => n9423, QN => n377);
   REGISTERS_reg_9_21_inst : DFFR_X1 port map( D => n6615, CK => CLK, RN => 
                           n3235, Q => n9424, QN => n378);
   REGISTERS_reg_9_20_inst : DFFR_X1 port map( D => n6616, CK => CLK, RN => 
                           n3235, Q => n9425, QN => n379);
   REGISTERS_reg_9_19_inst : DFFR_X1 port map( D => n6617, CK => CLK, RN => 
                           n3235, Q => n9426, QN => n380);
   REGISTERS_reg_9_18_inst : DFFR_X1 port map( D => n6618, CK => CLK, RN => 
                           n3235, Q => n9427, QN => n381);
   REGISTERS_reg_9_17_inst : DFFR_X1 port map( D => n6619, CK => CLK, RN => 
                           n3235, Q => n9428, QN => n382);
   REGISTERS_reg_9_16_inst : DFFR_X1 port map( D => n6620, CK => CLK, RN => 
                           n3235, Q => n9429, QN => n383);
   REGISTERS_reg_9_15_inst : DFFR_X1 port map( D => n6621, CK => CLK, RN => 
                           n3233, Q => n9430, QN => n384);
   REGISTERS_reg_9_14_inst : DFFR_X1 port map( D => n6622, CK => CLK, RN => 
                           n3233, Q => n9431, QN => n385);
   REGISTERS_reg_9_13_inst : DFFR_X1 port map( D => n6623, CK => CLK, RN => 
                           n3233, Q => n9432, QN => n386);
   REGISTERS_reg_9_12_inst : DFFR_X1 port map( D => n6624, CK => CLK, RN => 
                           n3233, Q => n9433, QN => n387);
   REGISTERS_reg_9_11_inst : DFFR_X1 port map( D => n6625, CK => CLK, RN => 
                           n3233, Q => n9434, QN => n388);
   REGISTERS_reg_9_10_inst : DFFR_X1 port map( D => n6626, CK => CLK, RN => 
                           n3233, Q => n9435, QN => n389);
   REGISTERS_reg_9_9_inst : DFFR_X1 port map( D => n6627, CK => CLK, RN => 
                           n3233, Q => n9436, QN => n390);
   REGISTERS_reg_9_8_inst : DFFR_X1 port map( D => n6628, CK => CLK, RN => 
                           n3233, Q => n9437, QN => n391);
   REGISTERS_reg_9_7_inst : DFFR_X1 port map( D => n6629, CK => CLK, RN => 
                           n3233, Q => n9438, QN => n392);
   REGISTERS_reg_9_6_inst : DFFR_X1 port map( D => n6630, CK => CLK, RN => 
                           n3233, Q => n9439, QN => n393);
   REGISTERS_reg_9_5_inst : DFFR_X1 port map( D => n6631, CK => CLK, RN => 
                           n3233, Q => n9440, QN => n394);
   REGISTERS_reg_9_4_inst : DFFR_X1 port map( D => n6632, CK => CLK, RN => 
                           n3233, Q => n9441, QN => n395);
   REGISTERS_reg_9_3_inst : DFFR_X1 port map( D => n6633, CK => CLK, RN => 
                           n3232, Q => n9442, QN => n396);
   REGISTERS_reg_9_2_inst : DFFR_X1 port map( D => n6634, CK => CLK, RN => 
                           n3232, Q => n9443, QN => n397);
   REGISTERS_reg_9_1_inst : DFFR_X1 port map( D => n6635, CK => CLK, RN => 
                           n3232, Q => n9444, QN => n398);
   REGISTERS_reg_9_0_inst : DFFR_X1 port map( D => n6636, CK => CLK, RN => 
                           n3232, Q => n9445, QN => n399);
   REGISTERS_reg_10_31_inst : DFFR_X1 port map( D => n6637, CK => CLK, RN => 
                           n3232, Q => n9446, QN => n400);
   REGISTERS_reg_10_30_inst : DFFR_X1 port map( D => n6638, CK => CLK, RN => 
                           n3232, Q => n9447, QN => n401);
   REGISTERS_reg_10_29_inst : DFFR_X1 port map( D => n6639, CK => CLK, RN => 
                           n3232, Q => n9448, QN => n402);
   REGISTERS_reg_10_28_inst : DFFR_X1 port map( D => n6640, CK => CLK, RN => 
                           n3232, Q => n9449, QN => n403);
   REGISTERS_reg_10_27_inst : DFFR_X1 port map( D => n6641, CK => CLK, RN => 
                           n3232, Q => n9450, QN => n404);
   REGISTERS_reg_10_26_inst : DFFR_X1 port map( D => n6642, CK => CLK, RN => 
                           n3232, Q => n9451, QN => n405);
   REGISTERS_reg_10_25_inst : DFFR_X1 port map( D => n6643, CK => CLK, RN => 
                           n3232, Q => n9452, QN => n406);
   REGISTERS_reg_10_24_inst : DFFR_X1 port map( D => n6644, CK => CLK, RN => 
                           n3232, Q => n9453, QN => n407);
   REGISTERS_reg_10_23_inst : DFFR_X1 port map( D => n6645, CK => CLK, RN => 
                           n3231, Q => n9454, QN => n408);
   REGISTERS_reg_10_22_inst : DFFR_X1 port map( D => n6646, CK => CLK, RN => 
                           n3231, Q => n9455, QN => n409);
   REGISTERS_reg_10_21_inst : DFFR_X1 port map( D => n6647, CK => CLK, RN => 
                           n3231, Q => n9456, QN => n410);
   REGISTERS_reg_10_20_inst : DFFR_X1 port map( D => n6648, CK => CLK, RN => 
                           n3231, Q => n9457, QN => n411);
   REGISTERS_reg_10_19_inst : DFFR_X1 port map( D => n6649, CK => CLK, RN => 
                           n3231, Q => n9458, QN => n412);
   REGISTERS_reg_10_18_inst : DFFR_X1 port map( D => n6650, CK => CLK, RN => 
                           n3231, Q => n9459, QN => n413);
   REGISTERS_reg_10_17_inst : DFFR_X1 port map( D => n6651, CK => CLK, RN => 
                           n3231, Q => n9460, QN => n414);
   REGISTERS_reg_10_16_inst : DFFR_X1 port map( D => n6652, CK => CLK, RN => 
                           n3231, Q => n9461, QN => n415);
   REGISTERS_reg_10_15_inst : DFFR_X1 port map( D => n6653, CK => CLK, RN => 
                           n3231, Q => n9462, QN => n416);
   REGISTERS_reg_10_14_inst : DFFR_X1 port map( D => n6654, CK => CLK, RN => 
                           n3231, Q => n9463, QN => n417);
   REGISTERS_reg_10_13_inst : DFFR_X1 port map( D => n6655, CK => CLK, RN => 
                           n3231, Q => n9464, QN => n418);
   REGISTERS_reg_10_12_inst : DFFR_X1 port map( D => n6656, CK => CLK, RN => 
                           n3231, Q => n9465, QN => n419);
   REGISTERS_reg_10_11_inst : DFFR_X1 port map( D => n6657, CK => CLK, RN => 
                           n3229, Q => n9466, QN => n420);
   REGISTERS_reg_10_10_inst : DFFR_X1 port map( D => n6658, CK => CLK, RN => 
                           n3229, Q => n9467, QN => n421);
   REGISTERS_reg_10_9_inst : DFFR_X1 port map( D => n6659, CK => CLK, RN => 
                           n3229, Q => n9468, QN => n422);
   REGISTERS_reg_10_8_inst : DFFR_X1 port map( D => n6660, CK => CLK, RN => 
                           n3229, Q => n9469, QN => n423);
   REGISTERS_reg_10_7_inst : DFFR_X1 port map( D => n6661, CK => CLK, RN => 
                           n3229, Q => n9470, QN => n424);
   REGISTERS_reg_10_6_inst : DFFR_X1 port map( D => n6662, CK => CLK, RN => 
                           n3229, Q => n9471, QN => n425);
   REGISTERS_reg_10_5_inst : DFFR_X1 port map( D => n6663, CK => CLK, RN => 
                           n3229, Q => n9472, QN => n426);
   REGISTERS_reg_10_4_inst : DFFR_X1 port map( D => n6664, CK => CLK, RN => 
                           n3229, Q => n9473, QN => n427);
   REGISTERS_reg_10_3_inst : DFFR_X1 port map( D => n6665, CK => CLK, RN => 
                           n3229, Q => n9474, QN => n428);
   REGISTERS_reg_10_2_inst : DFFR_X1 port map( D => n6666, CK => CLK, RN => 
                           n3229, Q => n9475, QN => n429);
   REGISTERS_reg_10_1_inst : DFFR_X1 port map( D => n6667, CK => CLK, RN => 
                           n3229, Q => n9476, QN => n430);
   REGISTERS_reg_10_0_inst : DFFR_X1 port map( D => n6668, CK => CLK, RN => 
                           n3229, Q => n9477, QN => n431);
   REGISTERS_reg_13_31_inst : DFFR_X1 port map( D => n6733, CK => CLK, RN => 
                           n3221, Q => n9478, QN => n496);
   REGISTERS_reg_13_30_inst : DFFR_X1 port map( D => n6734, CK => CLK, RN => 
                           n3221, Q => n9479, QN => n497);
   REGISTERS_reg_13_29_inst : DFFR_X1 port map( D => n6735, CK => CLK, RN => 
                           n3221, Q => n9480, QN => n498);
   REGISTERS_reg_13_28_inst : DFFR_X1 port map( D => n6736, CK => CLK, RN => 
                           n3221, Q => n9481, QN => n499);
   REGISTERS_reg_13_27_inst : DFFR_X1 port map( D => n6737, CK => CLK, RN => 
                           n3221, Q => n9482, QN => n500);
   REGISTERS_reg_13_26_inst : DFFR_X1 port map( D => n6738, CK => CLK, RN => 
                           n3221, Q => n9483, QN => n501);
   REGISTERS_reg_13_25_inst : DFFR_X1 port map( D => n6739, CK => CLK, RN => 
                           n3221, Q => n9484, QN => n502);
   REGISTERS_reg_13_24_inst : DFFR_X1 port map( D => n6740, CK => CLK, RN => 
                           n3221, Q => n9485, QN => n503);
   REGISTERS_reg_13_23_inst : DFFR_X1 port map( D => n6741, CK => CLK, RN => 
                           n3220, Q => n9486, QN => n504);
   REGISTERS_reg_13_22_inst : DFFR_X1 port map( D => n6742, CK => CLK, RN => 
                           n3220, Q => n9487, QN => n505);
   REGISTERS_reg_13_21_inst : DFFR_X1 port map( D => n6743, CK => CLK, RN => 
                           n3220, Q => n9488, QN => n506);
   REGISTERS_reg_13_20_inst : DFFR_X1 port map( D => n6744, CK => CLK, RN => 
                           n3220, Q => n9489, QN => n507);
   REGISTERS_reg_13_19_inst : DFFR_X1 port map( D => n6745, CK => CLK, RN => 
                           n3220, Q => n9490, QN => n508);
   REGISTERS_reg_13_18_inst : DFFR_X1 port map( D => n6746, CK => CLK, RN => 
                           n3220, Q => n9491, QN => n509);
   REGISTERS_reg_13_17_inst : DFFR_X1 port map( D => n6747, CK => CLK, RN => 
                           n3220, Q => n9492, QN => n510);
   REGISTERS_reg_13_16_inst : DFFR_X1 port map( D => n6748, CK => CLK, RN => 
                           n3220, Q => n9493, QN => n511);
   REGISTERS_reg_13_15_inst : DFFR_X1 port map( D => n6749, CK => CLK, RN => 
                           n3220, Q => n9494, QN => n512);
   REGISTERS_reg_13_14_inst : DFFR_X1 port map( D => n6750, CK => CLK, RN => 
                           n3220, Q => n9495, QN => n513);
   REGISTERS_reg_13_13_inst : DFFR_X1 port map( D => n6751, CK => CLK, RN => 
                           n3220, Q => n9496, QN => n514);
   REGISTERS_reg_13_12_inst : DFFR_X1 port map( D => n6752, CK => CLK, RN => 
                           n3220, Q => n9497, QN => n515);
   REGISTERS_reg_13_11_inst : DFFR_X1 port map( D => n6753, CK => CLK, RN => 
                           n3219, Q => n9498, QN => n516);
   REGISTERS_reg_13_10_inst : DFFR_X1 port map( D => n6754, CK => CLK, RN => 
                           n3219, Q => n9499, QN => n517);
   REGISTERS_reg_13_9_inst : DFFR_X1 port map( D => n6755, CK => CLK, RN => 
                           n3219, Q => n9500, QN => n518);
   REGISTERS_reg_13_8_inst : DFFR_X1 port map( D => n6756, CK => CLK, RN => 
                           n3219, Q => n9501, QN => n519);
   REGISTERS_reg_13_7_inst : DFFR_X1 port map( D => n6757, CK => CLK, RN => 
                           n3219, Q => n9502, QN => n520);
   REGISTERS_reg_13_6_inst : DFFR_X1 port map( D => n6758, CK => CLK, RN => 
                           n3219, Q => n9503, QN => n521);
   REGISTERS_reg_13_5_inst : DFFR_X1 port map( D => n6759, CK => CLK, RN => 
                           n3219, Q => n9504, QN => n522);
   REGISTERS_reg_13_4_inst : DFFR_X1 port map( D => n6760, CK => CLK, RN => 
                           n3219, Q => n9505, QN => n523);
   REGISTERS_reg_13_3_inst : DFFR_X1 port map( D => n6761, CK => CLK, RN => 
                           n3219, Q => n9506, QN => n524);
   REGISTERS_reg_13_2_inst : DFFR_X1 port map( D => n6762, CK => CLK, RN => 
                           n3219, Q => n9507, QN => n525);
   REGISTERS_reg_13_1_inst : DFFR_X1 port map( D => n6763, CK => CLK, RN => 
                           n3219, Q => n9508, QN => n526);
   REGISTERS_reg_13_0_inst : DFFR_X1 port map( D => n6764, CK => CLK, RN => 
                           n3219, Q => n9509, QN => n527);
   REGISTERS_reg_14_31_inst : DFFR_X1 port map( D => n6765, CK => CLK, RN => 
                           n3217, Q => n9510, QN => n528);
   REGISTERS_reg_14_30_inst : DFFR_X1 port map( D => n6766, CK => CLK, RN => 
                           n3217, Q => n9511, QN => n529);
   REGISTERS_reg_14_29_inst : DFFR_X1 port map( D => n6767, CK => CLK, RN => 
                           n3217, Q => n9512, QN => n530);
   REGISTERS_reg_14_28_inst : DFFR_X1 port map( D => n6768, CK => CLK, RN => 
                           n3217, Q => n9513, QN => n531);
   REGISTERS_reg_14_27_inst : DFFR_X1 port map( D => n6769, CK => CLK, RN => 
                           n3217, Q => n9514, QN => n532);
   REGISTERS_reg_14_26_inst : DFFR_X1 port map( D => n6770, CK => CLK, RN => 
                           n3217, Q => n9515, QN => n533);
   REGISTERS_reg_14_25_inst : DFFR_X1 port map( D => n6771, CK => CLK, RN => 
                           n3217, Q => n9516, QN => n534);
   REGISTERS_reg_14_24_inst : DFFR_X1 port map( D => n6772, CK => CLK, RN => 
                           n3217, Q => n9517, QN => n535);
   REGISTERS_reg_14_23_inst : DFFR_X1 port map( D => n6773, CK => CLK, RN => 
                           n3217, Q => n9518, QN => n536);
   REGISTERS_reg_14_22_inst : DFFR_X1 port map( D => n6774, CK => CLK, RN => 
                           n3217, Q => n9519, QN => n537);
   REGISTERS_reg_14_21_inst : DFFR_X1 port map( D => n6775, CK => CLK, RN => 
                           n3217, Q => n9520, QN => n538);
   REGISTERS_reg_14_20_inst : DFFR_X1 port map( D => n6776, CK => CLK, RN => 
                           n3217, Q => n9521, QN => n539);
   REGISTERS_reg_14_19_inst : DFFR_X1 port map( D => n6777, CK => CLK, RN => 
                           n3216, Q => n9522, QN => n540);
   REGISTERS_reg_14_18_inst : DFFR_X1 port map( D => n6778, CK => CLK, RN => 
                           n3216, Q => n9523, QN => n541);
   REGISTERS_reg_14_17_inst : DFFR_X1 port map( D => n6779, CK => CLK, RN => 
                           n3216, Q => n9524, QN => n542);
   REGISTERS_reg_14_16_inst : DFFR_X1 port map( D => n6780, CK => CLK, RN => 
                           n3216, Q => n9525, QN => n543);
   REGISTERS_reg_14_15_inst : DFFR_X1 port map( D => n6781, CK => CLK, RN => 
                           n3216, Q => n9526, QN => n544);
   REGISTERS_reg_14_14_inst : DFFR_X1 port map( D => n6782, CK => CLK, RN => 
                           n3216, Q => n9527, QN => n545);
   REGISTERS_reg_14_13_inst : DFFR_X1 port map( D => n6783, CK => CLK, RN => 
                           n3216, Q => n9528, QN => n546);
   REGISTERS_reg_14_12_inst : DFFR_X1 port map( D => n6784, CK => CLK, RN => 
                           n3216, Q => n9529, QN => n547);
   REGISTERS_reg_14_11_inst : DFFR_X1 port map( D => n6785, CK => CLK, RN => 
                           n3216, Q => n9530, QN => n548);
   REGISTERS_reg_14_10_inst : DFFR_X1 port map( D => n6786, CK => CLK, RN => 
                           n3216, Q => n9531, QN => n549);
   REGISTERS_reg_14_9_inst : DFFR_X1 port map( D => n6787, CK => CLK, RN => 
                           n3216, Q => n9532, QN => n550);
   REGISTERS_reg_14_8_inst : DFFR_X1 port map( D => n6788, CK => CLK, RN => 
                           n3216, Q => n9533, QN => n551);
   REGISTERS_reg_14_7_inst : DFFR_X1 port map( D => n6789, CK => CLK, RN => 
                           n3215, Q => n9534, QN => n552);
   REGISTERS_reg_14_6_inst : DFFR_X1 port map( D => n6790, CK => CLK, RN => 
                           n3215, Q => n9535, QN => n553);
   REGISTERS_reg_14_5_inst : DFFR_X1 port map( D => n6791, CK => CLK, RN => 
                           n3215, Q => n9536, QN => n554);
   REGISTERS_reg_14_4_inst : DFFR_X1 port map( D => n6792, CK => CLK, RN => 
                           n3215, Q => n9537, QN => n555);
   REGISTERS_reg_14_3_inst : DFFR_X1 port map( D => n6793, CK => CLK, RN => 
                           n3215, Q => n9538, QN => n556);
   REGISTERS_reg_14_2_inst : DFFR_X1 port map( D => n6794, CK => CLK, RN => 
                           n3215, Q => n9539, QN => n557);
   REGISTERS_reg_14_1_inst : DFFR_X1 port map( D => n6795, CK => CLK, RN => 
                           n3215, Q => n9540, QN => n558);
   REGISTERS_reg_14_0_inst : DFFR_X1 port map( D => n6796, CK => CLK, RN => 
                           n3215, Q => n9541, QN => n559);
   REGISTERS_reg_15_31_inst : DFFR_X1 port map( D => n6797, CK => CLK, RN => 
                           n3215, Q => n9542, QN => n560);
   REGISTERS_reg_15_30_inst : DFFR_X1 port map( D => n6798, CK => CLK, RN => 
                           n3215, Q => n9543, QN => n561);
   REGISTERS_reg_15_29_inst : DFFR_X1 port map( D => n6799, CK => CLK, RN => 
                           n3215, Q => n9544, QN => n562);
   REGISTERS_reg_15_28_inst : DFFR_X1 port map( D => n6800, CK => CLK, RN => 
                           n3215, Q => n9545, QN => n563);
   REGISTERS_reg_15_27_inst : DFFR_X1 port map( D => n6801, CK => CLK, RN => 
                           n3213, Q => n9546, QN => n564);
   REGISTERS_reg_15_26_inst : DFFR_X1 port map( D => n6802, CK => CLK, RN => 
                           n3213, Q => n9547, QN => n565);
   REGISTERS_reg_15_25_inst : DFFR_X1 port map( D => n6803, CK => CLK, RN => 
                           n3213, Q => n9548, QN => n566);
   REGISTERS_reg_15_24_inst : DFFR_X1 port map( D => n6804, CK => CLK, RN => 
                           n3213, Q => n9549, QN => n567);
   REGISTERS_reg_15_23_inst : DFFR_X1 port map( D => n6805, CK => CLK, RN => 
                           n3213, Q => n9550, QN => n568);
   REGISTERS_reg_15_22_inst : DFFR_X1 port map( D => n6806, CK => CLK, RN => 
                           n3213, Q => n9551, QN => n569);
   REGISTERS_reg_15_21_inst : DFFR_X1 port map( D => n6807, CK => CLK, RN => 
                           n3213, Q => n9552, QN => n570);
   REGISTERS_reg_15_20_inst : DFFR_X1 port map( D => n6808, CK => CLK, RN => 
                           n3213, Q => n9553, QN => n571);
   REGISTERS_reg_15_19_inst : DFFR_X1 port map( D => n6809, CK => CLK, RN => 
                           n3213, Q => n9554, QN => n572);
   REGISTERS_reg_15_18_inst : DFFR_X1 port map( D => n6810, CK => CLK, RN => 
                           n3213, Q => n9555, QN => n573);
   REGISTERS_reg_15_17_inst : DFFR_X1 port map( D => n6811, CK => CLK, RN => 
                           n3213, Q => n9556, QN => n574);
   REGISTERS_reg_15_16_inst : DFFR_X1 port map( D => n6812, CK => CLK, RN => 
                           n3213, Q => n9557, QN => n575);
   REGISTERS_reg_15_15_inst : DFFR_X1 port map( D => n6813, CK => CLK, RN => 
                           n3212, Q => n9558, QN => n576);
   REGISTERS_reg_15_14_inst : DFFR_X1 port map( D => n6814, CK => CLK, RN => 
                           n3212, Q => n9559, QN => n577);
   REGISTERS_reg_15_13_inst : DFFR_X1 port map( D => n6815, CK => CLK, RN => 
                           n3212, Q => n9560, QN => n578);
   REGISTERS_reg_15_12_inst : DFFR_X1 port map( D => n6816, CK => CLK, RN => 
                           n3212, Q => n9561, QN => n579);
   REGISTERS_reg_15_11_inst : DFFR_X1 port map( D => n6817, CK => CLK, RN => 
                           n3212, Q => n9562, QN => n580);
   REGISTERS_reg_15_10_inst : DFFR_X1 port map( D => n6818, CK => CLK, RN => 
                           n3212, Q => n9563, QN => n581);
   REGISTERS_reg_15_9_inst : DFFR_X1 port map( D => n6819, CK => CLK, RN => 
                           n3212, Q => n9564, QN => n582);
   REGISTERS_reg_15_8_inst : DFFR_X1 port map( D => n6820, CK => CLK, RN => 
                           n3212, Q => n9565, QN => n583);
   REGISTERS_reg_15_7_inst : DFFR_X1 port map( D => n6821, CK => CLK, RN => 
                           n3212, Q => n9566, QN => n584);
   REGISTERS_reg_15_6_inst : DFFR_X1 port map( D => n6822, CK => CLK, RN => 
                           n3212, Q => n9567, QN => n585);
   REGISTERS_reg_15_5_inst : DFFR_X1 port map( D => n6823, CK => CLK, RN => 
                           n3212, Q => n9568, QN => n586);
   REGISTERS_reg_15_4_inst : DFFR_X1 port map( D => n6824, CK => CLK, RN => 
                           n3212, Q => n9569, QN => n587);
   REGISTERS_reg_15_3_inst : DFFR_X1 port map( D => n6825, CK => CLK, RN => 
                           n3211, Q => n9570, QN => n588);
   REGISTERS_reg_15_2_inst : DFFR_X1 port map( D => n6826, CK => CLK, RN => 
                           n3211, Q => n9571, QN => n589);
   REGISTERS_reg_15_1_inst : DFFR_X1 port map( D => n6827, CK => CLK, RN => 
                           n3211, Q => n9572, QN => n590);
   REGISTERS_reg_15_0_inst : DFFR_X1 port map( D => n6828, CK => CLK, RN => 
                           n3211, Q => n9573, QN => n591);
   REGISTERS_reg_22_31_inst : DFFR_X1 port map( D => n7021, CK => CLK, RN => 
                           n3189, Q => n9574, QN => n784);
   REGISTERS_reg_22_30_inst : DFFR_X1 port map( D => n7022, CK => CLK, RN => 
                           n3189, Q => n9575, QN => n785);
   REGISTERS_reg_22_29_inst : DFFR_X1 port map( D => n7023, CK => CLK, RN => 
                           n3189, Q => n9576, QN => n786);
   REGISTERS_reg_22_28_inst : DFFR_X1 port map( D => n7024, CK => CLK, RN => 
                           n3189, Q => n9577, QN => n787);
   REGISTERS_reg_22_27_inst : DFFR_X1 port map( D => n7025, CK => CLK, RN => 
                           n3189, Q => n9578, QN => n788);
   REGISTERS_reg_22_26_inst : DFFR_X1 port map( D => n7026, CK => CLK, RN => 
                           n3189, Q => n9579, QN => n789);
   REGISTERS_reg_22_25_inst : DFFR_X1 port map( D => n7027, CK => CLK, RN => 
                           n3189, Q => n9580, QN => n790);
   REGISTERS_reg_22_24_inst : DFFR_X1 port map( D => n7028, CK => CLK, RN => 
                           n3189, Q => n9581, QN => n791);
   REGISTERS_reg_22_23_inst : DFFR_X1 port map( D => n7029, CK => CLK, RN => 
                           n3188, Q => n9582, QN => n792);
   REGISTERS_reg_22_22_inst : DFFR_X1 port map( D => n7030, CK => CLK, RN => 
                           n3188, Q => n9583, QN => n793);
   REGISTERS_reg_22_21_inst : DFFR_X1 port map( D => n7031, CK => CLK, RN => 
                           n3188, Q => n9584, QN => n794);
   REGISTERS_reg_22_20_inst : DFFR_X1 port map( D => n7032, CK => CLK, RN => 
                           n3188, Q => n9585, QN => n795);
   REGISTERS_reg_22_19_inst : DFFR_X1 port map( D => n7033, CK => CLK, RN => 
                           n3188, Q => n9586, QN => n796);
   REGISTERS_reg_22_18_inst : DFFR_X1 port map( D => n7034, CK => CLK, RN => 
                           n3188, Q => n9587, QN => n797);
   REGISTERS_reg_22_17_inst : DFFR_X1 port map( D => n7035, CK => CLK, RN => 
                           n3188, Q => n9588, QN => n798);
   REGISTERS_reg_22_16_inst : DFFR_X1 port map( D => n7036, CK => CLK, RN => 
                           n3188, Q => n9589, QN => n799);
   REGISTERS_reg_22_15_inst : DFFR_X1 port map( D => n7037, CK => CLK, RN => 
                           n3188, Q => n9590, QN => n800);
   REGISTERS_reg_22_14_inst : DFFR_X1 port map( D => n7038, CK => CLK, RN => 
                           n3188, Q => n9591, QN => n801);
   REGISTERS_reg_22_13_inst : DFFR_X1 port map( D => n7039, CK => CLK, RN => 
                           n3188, Q => n9592, QN => n802);
   REGISTERS_reg_22_12_inst : DFFR_X1 port map( D => n7040, CK => CLK, RN => 
                           n3188, Q => n9593, QN => n803);
   REGISTERS_reg_22_11_inst : DFFR_X1 port map( D => n7041, CK => CLK, RN => 
                           n3187, Q => n9594, QN => n804);
   REGISTERS_reg_22_10_inst : DFFR_X1 port map( D => n7042, CK => CLK, RN => 
                           n3187, Q => n9595, QN => n805);
   REGISTERS_reg_22_9_inst : DFFR_X1 port map( D => n7043, CK => CLK, RN => 
                           n3187, Q => n9596, QN => n806);
   REGISTERS_reg_22_8_inst : DFFR_X1 port map( D => n7044, CK => CLK, RN => 
                           n3187, Q => n9597, QN => n807);
   REGISTERS_reg_22_7_inst : DFFR_X1 port map( D => n7045, CK => CLK, RN => 
                           n3187, Q => n9598, QN => n808);
   REGISTERS_reg_22_6_inst : DFFR_X1 port map( D => n7046, CK => CLK, RN => 
                           n3187, Q => n9599, QN => n809);
   REGISTERS_reg_22_5_inst : DFFR_X1 port map( D => n7047, CK => CLK, RN => 
                           n3187, Q => n9600, QN => n810);
   REGISTERS_reg_22_4_inst : DFFR_X1 port map( D => n7048, CK => CLK, RN => 
                           n3187, Q => n9601, QN => n811);
   REGISTERS_reg_22_3_inst : DFFR_X1 port map( D => n7049, CK => CLK, RN => 
                           n3187, Q => n9602, QN => n812);
   REGISTERS_reg_22_2_inst : DFFR_X1 port map( D => n7050, CK => CLK, RN => 
                           n3187, Q => n9603, QN => n813);
   REGISTERS_reg_22_1_inst : DFFR_X1 port map( D => n7051, CK => CLK, RN => 
                           n3187, Q => n9604, QN => n814);
   REGISTERS_reg_22_0_inst : DFFR_X1 port map( D => n7052, CK => CLK, RN => 
                           n3187, Q => n9605, QN => n815);
   REGISTERS_reg_23_31_inst : DFFR_X1 port map( D => n7053, CK => CLK, RN => 
                           n3185, Q => n9606, QN => n816);
   REGISTERS_reg_23_30_inst : DFFR_X1 port map( D => n7054, CK => CLK, RN => 
                           n3185, Q => n9607, QN => n817);
   REGISTERS_reg_23_29_inst : DFFR_X1 port map( D => n7055, CK => CLK, RN => 
                           n3185, Q => n9608, QN => n818);
   REGISTERS_reg_23_28_inst : DFFR_X1 port map( D => n7056, CK => CLK, RN => 
                           n3185, Q => n9609, QN => n819);
   REGISTERS_reg_23_27_inst : DFFR_X1 port map( D => n7057, CK => CLK, RN => 
                           n3185, Q => n9610, QN => n820);
   REGISTERS_reg_23_26_inst : DFFR_X1 port map( D => n7058, CK => CLK, RN => 
                           n3185, Q => n9611, QN => n821);
   REGISTERS_reg_23_25_inst : DFFR_X1 port map( D => n7059, CK => CLK, RN => 
                           n3185, Q => n9612, QN => n822);
   REGISTERS_reg_23_24_inst : DFFR_X1 port map( D => n7060, CK => CLK, RN => 
                           n3185, Q => n9613, QN => n823);
   REGISTERS_reg_23_23_inst : DFFR_X1 port map( D => n7061, CK => CLK, RN => 
                           n3185, Q => n9614, QN => n824);
   REGISTERS_reg_23_22_inst : DFFR_X1 port map( D => n7062, CK => CLK, RN => 
                           n3185, Q => n9615, QN => n825);
   REGISTERS_reg_23_21_inst : DFFR_X1 port map( D => n7063, CK => CLK, RN => 
                           n3185, Q => n9616, QN => n826);
   REGISTERS_reg_23_20_inst : DFFR_X1 port map( D => n7064, CK => CLK, RN => 
                           n3185, Q => n9617, QN => n827);
   REGISTERS_reg_23_19_inst : DFFR_X1 port map( D => n7065, CK => CLK, RN => 
                           n3184, Q => n9618, QN => n828);
   REGISTERS_reg_23_18_inst : DFFR_X1 port map( D => n7066, CK => CLK, RN => 
                           n3184, Q => n9619, QN => n829);
   REGISTERS_reg_23_17_inst : DFFR_X1 port map( D => n7067, CK => CLK, RN => 
                           n3184, Q => n9620, QN => n830);
   REGISTERS_reg_23_16_inst : DFFR_X1 port map( D => n7068, CK => CLK, RN => 
                           n3184, Q => n9621, QN => n831);
   REGISTERS_reg_23_15_inst : DFFR_X1 port map( D => n7069, CK => CLK, RN => 
                           n3184, Q => n9622, QN => n832);
   REGISTERS_reg_23_14_inst : DFFR_X1 port map( D => n7070, CK => CLK, RN => 
                           n3184, Q => n9623, QN => n833);
   REGISTERS_reg_23_13_inst : DFFR_X1 port map( D => n7071, CK => CLK, RN => 
                           n3184, Q => n9624, QN => n834);
   REGISTERS_reg_23_12_inst : DFFR_X1 port map( D => n7072, CK => CLK, RN => 
                           n3184, Q => n9625, QN => n835);
   REGISTERS_reg_23_11_inst : DFFR_X1 port map( D => n7073, CK => CLK, RN => 
                           n3184, Q => n9626, QN => n836);
   REGISTERS_reg_23_10_inst : DFFR_X1 port map( D => n7074, CK => CLK, RN => 
                           n3184, Q => n9627, QN => n837);
   REGISTERS_reg_23_9_inst : DFFR_X1 port map( D => n7075, CK => CLK, RN => 
                           n3184, Q => n9628, QN => n838);
   REGISTERS_reg_23_8_inst : DFFR_X1 port map( D => n7076, CK => CLK, RN => 
                           n3184, Q => n9629, QN => n839);
   REGISTERS_reg_23_7_inst : DFFR_X1 port map( D => n7077, CK => CLK, RN => 
                           n3183, Q => n9630, QN => n840);
   REGISTERS_reg_23_6_inst : DFFR_X1 port map( D => n7078, CK => CLK, RN => 
                           n3183, Q => n9631, QN => n841);
   REGISTERS_reg_23_5_inst : DFFR_X1 port map( D => n7079, CK => CLK, RN => 
                           n3183, Q => n9632, QN => n842);
   REGISTERS_reg_23_4_inst : DFFR_X1 port map( D => n7080, CK => CLK, RN => 
                           n3183, Q => n9633, QN => n843);
   REGISTERS_reg_23_3_inst : DFFR_X1 port map( D => n7081, CK => CLK, RN => 
                           n3183, Q => n9634, QN => n844);
   REGISTERS_reg_23_2_inst : DFFR_X1 port map( D => n7082, CK => CLK, RN => 
                           n3183, Q => n9635, QN => n845);
   REGISTERS_reg_23_1_inst : DFFR_X1 port map( D => n7083, CK => CLK, RN => 
                           n3183, Q => n9636, QN => n846);
   REGISTERS_reg_23_0_inst : DFFR_X1 port map( D => n7084, CK => CLK, RN => 
                           n3183, Q => n9637, QN => n847);
   REGISTERS_reg_24_31_inst : DFFR_X1 port map( D => n7085, CK => CLK, RN => 
                           n3183, Q => n9638, QN => n848);
   REGISTERS_reg_24_30_inst : DFFR_X1 port map( D => n7086, CK => CLK, RN => 
                           n3183, Q => n9639, QN => n849);
   REGISTERS_reg_24_29_inst : DFFR_X1 port map( D => n7087, CK => CLK, RN => 
                           n3183, Q => n9640, QN => n850);
   REGISTERS_reg_24_28_inst : DFFR_X1 port map( D => n7088, CK => CLK, RN => 
                           n3183, Q => n9641, QN => n851);
   REGISTERS_reg_24_27_inst : DFFR_X1 port map( D => n7089, CK => CLK, RN => 
                           n3181, Q => n9642, QN => n852);
   REGISTERS_reg_24_26_inst : DFFR_X1 port map( D => n7090, CK => CLK, RN => 
                           n3181, Q => n9643, QN => n853);
   REGISTERS_reg_24_25_inst : DFFR_X1 port map( D => n7091, CK => CLK, RN => 
                           n3181, Q => n9644, QN => n854);
   REGISTERS_reg_24_24_inst : DFFR_X1 port map( D => n7092, CK => CLK, RN => 
                           n3181, Q => n9645, QN => n855);
   REGISTERS_reg_24_23_inst : DFFR_X1 port map( D => n7093, CK => CLK, RN => 
                           n3181, Q => n9646, QN => n856);
   REGISTERS_reg_24_22_inst : DFFR_X1 port map( D => n7094, CK => CLK, RN => 
                           n3181, Q => n9647, QN => n857);
   REGISTERS_reg_24_21_inst : DFFR_X1 port map( D => n7095, CK => CLK, RN => 
                           n3181, Q => n9648, QN => n858);
   REGISTERS_reg_24_20_inst : DFFR_X1 port map( D => n7096, CK => CLK, RN => 
                           n3181, Q => n9649, QN => n859);
   REGISTERS_reg_24_19_inst : DFFR_X1 port map( D => n7097, CK => CLK, RN => 
                           n3181, Q => n9650, QN => n860);
   REGISTERS_reg_24_18_inst : DFFR_X1 port map( D => n7098, CK => CLK, RN => 
                           n3181, Q => n9651, QN => n861);
   REGISTERS_reg_24_17_inst : DFFR_X1 port map( D => n7099, CK => CLK, RN => 
                           n3181, Q => n9652, QN => n862);
   REGISTERS_reg_24_16_inst : DFFR_X1 port map( D => n7100, CK => CLK, RN => 
                           n3181, Q => n9653, QN => n863);
   REGISTERS_reg_24_15_inst : DFFR_X1 port map( D => n7101, CK => CLK, RN => 
                           n3180, Q => n9654, QN => n864);
   REGISTERS_reg_24_14_inst : DFFR_X1 port map( D => n7102, CK => CLK, RN => 
                           n3180, Q => n9655, QN => n865);
   REGISTERS_reg_24_13_inst : DFFR_X1 port map( D => n7103, CK => CLK, RN => 
                           n3180, Q => n9656, QN => n866);
   REGISTERS_reg_24_12_inst : DFFR_X1 port map( D => n7104, CK => CLK, RN => 
                           n3180, Q => n9657, QN => n867);
   REGISTERS_reg_24_11_inst : DFFR_X1 port map( D => n7105, CK => CLK, RN => 
                           n3180, Q => n9658, QN => n868);
   REGISTERS_reg_24_10_inst : DFFR_X1 port map( D => n7106, CK => CLK, RN => 
                           n3180, Q => n9659, QN => n869);
   REGISTERS_reg_24_9_inst : DFFR_X1 port map( D => n7107, CK => CLK, RN => 
                           n3180, Q => n9660, QN => n870);
   REGISTERS_reg_24_8_inst : DFFR_X1 port map( D => n7108, CK => CLK, RN => 
                           n3180, Q => n9661, QN => n871);
   REGISTERS_reg_24_7_inst : DFFR_X1 port map( D => n7109, CK => CLK, RN => 
                           n3180, Q => n9662, QN => n872);
   REGISTERS_reg_24_6_inst : DFFR_X1 port map( D => n7110, CK => CLK, RN => 
                           n3180, Q => n9663, QN => n873);
   REGISTERS_reg_24_5_inst : DFFR_X1 port map( D => n7111, CK => CLK, RN => 
                           n3180, Q => n9664, QN => n874);
   REGISTERS_reg_24_4_inst : DFFR_X1 port map( D => n7112, CK => CLK, RN => 
                           n3180, Q => n9665, QN => n875);
   REGISTERS_reg_24_3_inst : DFFR_X1 port map( D => n7113, CK => CLK, RN => 
                           n3178, Q => n9666, QN => n876);
   REGISTERS_reg_24_2_inst : DFFR_X1 port map( D => n7114, CK => CLK, RN => 
                           n3178, Q => n9667, QN => n877);
   REGISTERS_reg_24_1_inst : DFFR_X1 port map( D => n7115, CK => CLK, RN => 
                           n3178, Q => n9668, QN => n878);
   REGISTERS_reg_24_0_inst : DFFR_X1 port map( D => n7116, CK => CLK, RN => 
                           n3178, Q => n9669, QN => n879);
   REGISTERS_reg_25_31_inst : DFFR_X1 port map( D => n7117, CK => CLK, RN => 
                           n3178, Q => n9670, QN => n880);
   REGISTERS_reg_25_30_inst : DFFR_X1 port map( D => n7118, CK => CLK, RN => 
                           n3178, Q => n9671, QN => n881);
   REGISTERS_reg_25_29_inst : DFFR_X1 port map( D => n7119, CK => CLK, RN => 
                           n3178, Q => n9672, QN => n882);
   REGISTERS_reg_25_28_inst : DFFR_X1 port map( D => n7120, CK => CLK, RN => 
                           n3178, Q => n9673, QN => n883);
   REGISTERS_reg_25_27_inst : DFFR_X1 port map( D => n7121, CK => CLK, RN => 
                           n3178, Q => n9674, QN => n884);
   REGISTERS_reg_25_26_inst : DFFR_X1 port map( D => n7122, CK => CLK, RN => 
                           n3178, Q => n9675, QN => n885);
   REGISTERS_reg_25_25_inst : DFFR_X1 port map( D => n7123, CK => CLK, RN => 
                           n3178, Q => n9676, QN => n886);
   REGISTERS_reg_25_24_inst : DFFR_X1 port map( D => n7124, CK => CLK, RN => 
                           n3178, Q => n9677, QN => n887);
   REGISTERS_reg_25_23_inst : DFFR_X1 port map( D => n7125, CK => CLK, RN => 
                           n3176, Q => n9678, QN => n888);
   REGISTERS_reg_25_22_inst : DFFR_X1 port map( D => n7126, CK => CLK, RN => 
                           n3176, Q => n9679, QN => n889);
   REGISTERS_reg_25_21_inst : DFFR_X1 port map( D => n7127, CK => CLK, RN => 
                           n3176, Q => n9680, QN => n890);
   REGISTERS_reg_25_20_inst : DFFR_X1 port map( D => n7128, CK => CLK, RN => 
                           n3176, Q => n9681, QN => n891);
   REGISTERS_reg_25_19_inst : DFFR_X1 port map( D => n7129, CK => CLK, RN => 
                           n3176, Q => n9682, QN => n892);
   REGISTERS_reg_25_18_inst : DFFR_X1 port map( D => n7130, CK => CLK, RN => 
                           n3176, Q => n9683, QN => n893);
   REGISTERS_reg_25_17_inst : DFFR_X1 port map( D => n7131, CK => CLK, RN => 
                           n3176, Q => n9684, QN => n894);
   REGISTERS_reg_25_16_inst : DFFR_X1 port map( D => n7132, CK => CLK, RN => 
                           n3176, Q => n9685, QN => n895);
   REGISTERS_reg_25_15_inst : DFFR_X1 port map( D => n7133, CK => CLK, RN => 
                           n3176, Q => n9686, QN => n896);
   REGISTERS_reg_25_14_inst : DFFR_X1 port map( D => n7134, CK => CLK, RN => 
                           n3176, Q => n9687, QN => n897);
   REGISTERS_reg_25_13_inst : DFFR_X1 port map( D => n7135, CK => CLK, RN => 
                           n3176, Q => n9688, QN => n898);
   REGISTERS_reg_25_12_inst : DFFR_X1 port map( D => n7136, CK => CLK, RN => 
                           n3176, Q => n9689, QN => n899);
   REGISTERS_reg_25_11_inst : DFFR_X1 port map( D => n7137, CK => CLK, RN => 
                           n3175, Q => n9690, QN => n900);
   REGISTERS_reg_25_10_inst : DFFR_X1 port map( D => n7138, CK => CLK, RN => 
                           n3175, Q => n9691, QN => n901);
   REGISTERS_reg_25_9_inst : DFFR_X1 port map( D => n7139, CK => CLK, RN => 
                           n3175, Q => n9692, QN => n902);
   REGISTERS_reg_25_8_inst : DFFR_X1 port map( D => n7140, CK => CLK, RN => 
                           n3175, Q => n9693, QN => n903);
   REGISTERS_reg_25_7_inst : DFFR_X1 port map( D => n7141, CK => CLK, RN => 
                           n3175, Q => n9694, QN => n904);
   REGISTERS_reg_25_6_inst : DFFR_X1 port map( D => n7142, CK => CLK, RN => 
                           n3175, Q => n9695, QN => n905);
   REGISTERS_reg_25_5_inst : DFFR_X1 port map( D => n7143, CK => CLK, RN => 
                           n3175, Q => n9696, QN => n906);
   REGISTERS_reg_25_4_inst : DFFR_X1 port map( D => n7144, CK => CLK, RN => 
                           n3175, Q => n9697, QN => n907);
   REGISTERS_reg_25_3_inst : DFFR_X1 port map( D => n7145, CK => CLK, RN => 
                           n3175, Q => n9698, QN => n908);
   REGISTERS_reg_25_2_inst : DFFR_X1 port map( D => n7146, CK => CLK, RN => 
                           n3175, Q => n9699, QN => n909);
   REGISTERS_reg_25_1_inst : DFFR_X1 port map( D => n7147, CK => CLK, RN => 
                           n3175, Q => n9700, QN => n910);
   REGISTERS_reg_25_0_inst : DFFR_X1 port map( D => n7148, CK => CLK, RN => 
                           n3175, Q => n9701, QN => n911);
   REGISTERS_reg_26_31_inst : DFFR_X1 port map( D => n7149, CK => CLK, RN => 
                           n3174, Q => n9702, QN => n912);
   REGISTERS_reg_26_30_inst : DFFR_X1 port map( D => n7150, CK => CLK, RN => 
                           n3174, Q => n9703, QN => n913);
   REGISTERS_reg_26_29_inst : DFFR_X1 port map( D => n7151, CK => CLK, RN => 
                           n3174, Q => n9704, QN => n914);
   REGISTERS_reg_26_28_inst : DFFR_X1 port map( D => n7152, CK => CLK, RN => 
                           n3174, Q => n9705, QN => n915);
   REGISTERS_reg_26_27_inst : DFFR_X1 port map( D => n7153, CK => CLK, RN => 
                           n3174, Q => n9706, QN => n916);
   REGISTERS_reg_26_26_inst : DFFR_X1 port map( D => n7154, CK => CLK, RN => 
                           n3174, Q => n9707, QN => n917);
   REGISTERS_reg_26_25_inst : DFFR_X1 port map( D => n7155, CK => CLK, RN => 
                           n3174, Q => n9708, QN => n918);
   REGISTERS_reg_26_24_inst : DFFR_X1 port map( D => n7156, CK => CLK, RN => 
                           n3174, Q => n9709, QN => n919);
   REGISTERS_reg_26_23_inst : DFFR_X1 port map( D => n7157, CK => CLK, RN => 
                           n3174, Q => n9710, QN => n920);
   REGISTERS_reg_26_22_inst : DFFR_X1 port map( D => n7158, CK => CLK, RN => 
                           n3174, Q => n9711, QN => n921);
   REGISTERS_reg_26_21_inst : DFFR_X1 port map( D => n7159, CK => CLK, RN => 
                           n3174, Q => n9712, QN => n922);
   REGISTERS_reg_26_20_inst : DFFR_X1 port map( D => n7160, CK => CLK, RN => 
                           n3174, Q => n9713, QN => n923);
   REGISTERS_reg_26_19_inst : DFFR_X1 port map( D => n7161, CK => CLK, RN => 
                           n3172, Q => n9714, QN => n924);
   REGISTERS_reg_26_18_inst : DFFR_X1 port map( D => n7162, CK => CLK, RN => 
                           n3172, Q => n9715, QN => n925);
   REGISTERS_reg_26_17_inst : DFFR_X1 port map( D => n7163, CK => CLK, RN => 
                           n3172, Q => n9716, QN => n926);
   REGISTERS_reg_26_16_inst : DFFR_X1 port map( D => n7164, CK => CLK, RN => 
                           n3172, Q => n9717, QN => n927);
   REGISTERS_reg_26_15_inst : DFFR_X1 port map( D => n7165, CK => CLK, RN => 
                           n3172, Q => n9718, QN => n928);
   REGISTERS_reg_26_14_inst : DFFR_X1 port map( D => n7166, CK => CLK, RN => 
                           n3172, Q => n9719, QN => n929);
   REGISTERS_reg_26_13_inst : DFFR_X1 port map( D => n7167, CK => CLK, RN => 
                           n3172, Q => n9720, QN => n930);
   REGISTERS_reg_26_12_inst : DFFR_X1 port map( D => n7168, CK => CLK, RN => 
                           n3172, Q => n9721, QN => n931);
   REGISTERS_reg_26_11_inst : DFFR_X1 port map( D => n7169, CK => CLK, RN => 
                           n3172, Q => n9722, QN => n932);
   REGISTERS_reg_26_10_inst : DFFR_X1 port map( D => n7170, CK => CLK, RN => 
                           n3172, Q => n9723, QN => n933);
   REGISTERS_reg_26_9_inst : DFFR_X1 port map( D => n7171, CK => CLK, RN => 
                           n3172, Q => n9724, QN => n934);
   REGISTERS_reg_26_8_inst : DFFR_X1 port map( D => n7172, CK => CLK, RN => 
                           n3172, Q => n9725, QN => n935);
   REGISTERS_reg_26_7_inst : DFFR_X1 port map( D => n7173, CK => CLK, RN => 
                           n3171, Q => n9726, QN => n936);
   REGISTERS_reg_26_6_inst : DFFR_X1 port map( D => n7174, CK => CLK, RN => 
                           n3171, Q => n9727, QN => n937);
   REGISTERS_reg_26_5_inst : DFFR_X1 port map( D => n7175, CK => CLK, RN => 
                           n3171, Q => n9728, QN => n938);
   REGISTERS_reg_26_4_inst : DFFR_X1 port map( D => n7176, CK => CLK, RN => 
                           n3171, Q => n9729, QN => n939);
   REGISTERS_reg_26_3_inst : DFFR_X1 port map( D => n7177, CK => CLK, RN => 
                           n3171, Q => n9730, QN => n940);
   REGISTERS_reg_26_2_inst : DFFR_X1 port map( D => n7178, CK => CLK, RN => 
                           n3171, Q => n9731, QN => n941);
   REGISTERS_reg_26_1_inst : DFFR_X1 port map( D => n7179, CK => CLK, RN => 
                           n3171, Q => n9732, QN => n942);
   REGISTERS_reg_26_0_inst : DFFR_X1 port map( D => n7180, CK => CLK, RN => 
                           n3171, Q => n9733, QN => n943);
   REGISTERS_reg_27_31_inst : DFFR_X1 port map( D => n7181, CK => CLK, RN => 
                           n3171, Q => n9734, QN => n944);
   REGISTERS_reg_27_30_inst : DFFR_X1 port map( D => n7182, CK => CLK, RN => 
                           n3171, Q => n9735, QN => n945);
   REGISTERS_reg_27_29_inst : DFFR_X1 port map( D => n7183, CK => CLK, RN => 
                           n3171, Q => n9736, QN => n946);
   REGISTERS_reg_27_28_inst : DFFR_X1 port map( D => n7184, CK => CLK, RN => 
                           n3171, Q => n9737, QN => n947);
   REGISTERS_reg_27_27_inst : DFFR_X1 port map( D => n7185, CK => CLK, RN => 
                           n3170, Q => n9738, QN => n948);
   REGISTERS_reg_27_26_inst : DFFR_X1 port map( D => n7186, CK => CLK, RN => 
                           n3170, Q => n9739, QN => n949);
   REGISTERS_reg_27_25_inst : DFFR_X1 port map( D => n7187, CK => CLK, RN => 
                           n3170, Q => n9740, QN => n950);
   REGISTERS_reg_27_24_inst : DFFR_X1 port map( D => n7188, CK => CLK, RN => 
                           n3170, Q => n9741, QN => n951);
   REGISTERS_reg_27_23_inst : DFFR_X1 port map( D => n7189, CK => CLK, RN => 
                           n3170, Q => n9742, QN => n952);
   REGISTERS_reg_27_22_inst : DFFR_X1 port map( D => n7190, CK => CLK, RN => 
                           n3170, Q => n9743, QN => n953);
   REGISTERS_reg_27_21_inst : DFFR_X1 port map( D => n7191, CK => CLK, RN => 
                           n3170, Q => n9744, QN => n954);
   REGISTERS_reg_27_20_inst : DFFR_X1 port map( D => n7192, CK => CLK, RN => 
                           n3170, Q => n9745, QN => n955);
   REGISTERS_reg_27_19_inst : DFFR_X1 port map( D => n7193, CK => CLK, RN => 
                           n3170, Q => n9746, QN => n956);
   REGISTERS_reg_27_18_inst : DFFR_X1 port map( D => n7194, CK => CLK, RN => 
                           n3170, Q => n9747, QN => n957);
   REGISTERS_reg_27_17_inst : DFFR_X1 port map( D => n7195, CK => CLK, RN => 
                           n3170, Q => n9748, QN => n958);
   REGISTERS_reg_27_16_inst : DFFR_X1 port map( D => n7196, CK => CLK, RN => 
                           n3170, Q => n9749, QN => n959);
   REGISTERS_reg_27_15_inst : DFFR_X1 port map( D => n7197, CK => CLK, RN => 
                           n3168, Q => n9750, QN => n960);
   REGISTERS_reg_27_14_inst : DFFR_X1 port map( D => n7198, CK => CLK, RN => 
                           n3168, Q => n9751, QN => n961);
   REGISTERS_reg_27_13_inst : DFFR_X1 port map( D => n7199, CK => CLK, RN => 
                           n3168, Q => n9752, QN => n962);
   REGISTERS_reg_27_12_inst : DFFR_X1 port map( D => n7200, CK => CLK, RN => 
                           n3168, Q => n9753, QN => n963);
   REGISTERS_reg_27_11_inst : DFFR_X1 port map( D => n7201, CK => CLK, RN => 
                           n3168, Q => n9754, QN => n964);
   REGISTERS_reg_27_10_inst : DFFR_X1 port map( D => n7202, CK => CLK, RN => 
                           n3168, Q => n9755, QN => n965);
   REGISTERS_reg_27_9_inst : DFFR_X1 port map( D => n7203, CK => CLK, RN => 
                           n3168, Q => n9756, QN => n966);
   REGISTERS_reg_27_8_inst : DFFR_X1 port map( D => n7204, CK => CLK, RN => 
                           n3168, Q => n9757, QN => n967);
   REGISTERS_reg_27_7_inst : DFFR_X1 port map( D => n7205, CK => CLK, RN => 
                           n3168, Q => n9758, QN => n968);
   REGISTERS_reg_27_6_inst : DFFR_X1 port map( D => n7206, CK => CLK, RN => 
                           n3168, Q => n9759, QN => n969);
   REGISTERS_reg_27_5_inst : DFFR_X1 port map( D => n7207, CK => CLK, RN => 
                           n3168, Q => n9760, QN => n970);
   REGISTERS_reg_27_4_inst : DFFR_X1 port map( D => n7208, CK => CLK, RN => 
                           n3168, Q => n9761, QN => n971);
   REGISTERS_reg_27_3_inst : DFFR_X1 port map( D => n7209, CK => CLK, RN => 
                           n3167, Q => n9762, QN => n972);
   REGISTERS_reg_27_2_inst : DFFR_X1 port map( D => n7210, CK => CLK, RN => 
                           n3167, Q => n9763, QN => n973);
   REGISTERS_reg_27_1_inst : DFFR_X1 port map( D => n7211, CK => CLK, RN => 
                           n3167, Q => n9764, QN => n974);
   REGISTERS_reg_27_0_inst : DFFR_X1 port map( D => n7212, CK => CLK, RN => 
                           n3167, Q => n9765, QN => n975);
   REGISTERS_reg_28_31_inst : DFFR_X1 port map( D => n7213, CK => CLK, RN => 
                           n3167, Q => n9766, QN => n976);
   REGISTERS_reg_28_30_inst : DFFR_X1 port map( D => n7214, CK => CLK, RN => 
                           n3167, Q => n9767, QN => n977);
   REGISTERS_reg_28_29_inst : DFFR_X1 port map( D => n7215, CK => CLK, RN => 
                           n3167, Q => n9768, QN => n978);
   REGISTERS_reg_28_28_inst : DFFR_X1 port map( D => n7216, CK => CLK, RN => 
                           n3167, Q => n9769, QN => n979);
   REGISTERS_reg_28_27_inst : DFFR_X1 port map( D => n7217, CK => CLK, RN => 
                           n3167, Q => n9770, QN => n980);
   REGISTERS_reg_28_26_inst : DFFR_X1 port map( D => n7218, CK => CLK, RN => 
                           n3167, Q => n9771, QN => n981);
   REGISTERS_reg_28_25_inst : DFFR_X1 port map( D => n7219, CK => CLK, RN => 
                           n3167, Q => n9772, QN => n982);
   REGISTERS_reg_28_24_inst : DFFR_X1 port map( D => n7220, CK => CLK, RN => 
                           n3167, Q => n9773, QN => n983);
   REGISTERS_reg_28_23_inst : DFFR_X1 port map( D => n7221, CK => CLK, RN => 
                           n3166, Q => n9774, QN => n984);
   REGISTERS_reg_28_22_inst : DFFR_X1 port map( D => n7222, CK => CLK, RN => 
                           n3166, Q => n9775, QN => n985);
   REGISTERS_reg_28_21_inst : DFFR_X1 port map( D => n7223, CK => CLK, RN => 
                           n3166, Q => n9776, QN => n986);
   REGISTERS_reg_28_20_inst : DFFR_X1 port map( D => n7224, CK => CLK, RN => 
                           n3166, Q => n9777, QN => n987);
   REGISTERS_reg_28_19_inst : DFFR_X1 port map( D => n7225, CK => CLK, RN => 
                           n3166, Q => n9778, QN => n988);
   REGISTERS_reg_28_18_inst : DFFR_X1 port map( D => n7226, CK => CLK, RN => 
                           n3166, Q => n9779, QN => n989);
   REGISTERS_reg_28_17_inst : DFFR_X1 port map( D => n7227, CK => CLK, RN => 
                           n3166, Q => n9780, QN => n990);
   REGISTERS_reg_28_16_inst : DFFR_X1 port map( D => n7228, CK => CLK, RN => 
                           n3166, Q => n9781, QN => n991);
   REGISTERS_reg_28_15_inst : DFFR_X1 port map( D => n7229, CK => CLK, RN => 
                           n3166, Q => n9782, QN => n992);
   REGISTERS_reg_28_14_inst : DFFR_X1 port map( D => n7230, CK => CLK, RN => 
                           n3166, Q => n9783, QN => n993);
   REGISTERS_reg_28_13_inst : DFFR_X1 port map( D => n7231, CK => CLK, RN => 
                           n3166, Q => n9784, QN => n994);
   REGISTERS_reg_28_12_inst : DFFR_X1 port map( D => n7232, CK => CLK, RN => 
                           n3166, Q => n9785, QN => n995);
   REGISTERS_reg_28_11_inst : DFFR_X1 port map( D => n7233, CK => CLK, RN => 
                           n3164, Q => n9786, QN => n996);
   REGISTERS_reg_28_10_inst : DFFR_X1 port map( D => n7234, CK => CLK, RN => 
                           n3164, Q => n9787, QN => n997);
   REGISTERS_reg_28_9_inst : DFFR_X1 port map( D => n7235, CK => CLK, RN => 
                           n3164, Q => n9788, QN => n998);
   REGISTERS_reg_28_8_inst : DFFR_X1 port map( D => n7236, CK => CLK, RN => 
                           n3164, Q => n9789, QN => n999);
   REGISTERS_reg_28_7_inst : DFFR_X1 port map( D => n7237, CK => CLK, RN => 
                           n3164, Q => n9790, QN => n1000);
   REGISTERS_reg_28_6_inst : DFFR_X1 port map( D => n7238, CK => CLK, RN => 
                           n3164, Q => n9791, QN => n1001);
   REGISTERS_reg_28_5_inst : DFFR_X1 port map( D => n7239, CK => CLK, RN => 
                           n3164, Q => n9792, QN => n1002);
   REGISTERS_reg_28_4_inst : DFFR_X1 port map( D => n7240, CK => CLK, RN => 
                           n3164, Q => n9793, QN => n1003);
   REGISTERS_reg_28_3_inst : DFFR_X1 port map( D => n7241, CK => CLK, RN => 
                           n3164, Q => n9794, QN => n1004);
   REGISTERS_reg_28_2_inst : DFFR_X1 port map( D => n7242, CK => CLK, RN => 
                           n3164, Q => n9795, QN => n1005);
   REGISTERS_reg_28_1_inst : DFFR_X1 port map( D => n7243, CK => CLK, RN => 
                           n3164, Q => n9796, QN => n1006);
   REGISTERS_reg_28_0_inst : DFFR_X1 port map( D => n7244, CK => CLK, RN => 
                           n3164, Q => n9797, QN => n1007);
   REGISTERS_reg_29_31_inst : DFFR_X1 port map( D => n7245, CK => CLK, RN => 
                           n3163, Q => n9798, QN => n1008);
   REGISTERS_reg_29_30_inst : DFFR_X1 port map( D => n7246, CK => CLK, RN => 
                           n3163, Q => n9799, QN => n1009);
   REGISTERS_reg_29_29_inst : DFFR_X1 port map( D => n7247, CK => CLK, RN => 
                           n3163, Q => n9800, QN => n1010);
   REGISTERS_reg_29_28_inst : DFFR_X1 port map( D => n7248, CK => CLK, RN => 
                           n3163, Q => n9801, QN => n1011);
   REGISTERS_reg_29_27_inst : DFFR_X1 port map( D => n7249, CK => CLK, RN => 
                           n3163, Q => n9802, QN => n1012);
   REGISTERS_reg_29_26_inst : DFFR_X1 port map( D => n7250, CK => CLK, RN => 
                           n3163, Q => n9803, QN => n1013);
   REGISTERS_reg_29_25_inst : DFFR_X1 port map( D => n7251, CK => CLK, RN => 
                           n3163, Q => n9804, QN => n1014);
   REGISTERS_reg_29_24_inst : DFFR_X1 port map( D => n7252, CK => CLK, RN => 
                           n3163, Q => n9805, QN => n1015);
   REGISTERS_reg_29_23_inst : DFFR_X1 port map( D => n7253, CK => CLK, RN => 
                           n3163, Q => n9806, QN => n1016);
   REGISTERS_reg_29_22_inst : DFFR_X1 port map( D => n7254, CK => CLK, RN => 
                           n3163, Q => n9807, QN => n1017);
   REGISTERS_reg_29_21_inst : DFFR_X1 port map( D => n7255, CK => CLK, RN => 
                           n3163, Q => n9808, QN => n1018);
   REGISTERS_reg_29_20_inst : DFFR_X1 port map( D => n7256, CK => CLK, RN => 
                           n3163, Q => n9809, QN => n1019);
   REGISTERS_reg_29_19_inst : DFFR_X1 port map( D => n7257, CK => CLK, RN => 
                           n3162, Q => n9810, QN => n1020);
   REGISTERS_reg_29_18_inst : DFFR_X1 port map( D => n7258, CK => CLK, RN => 
                           n3162, Q => n9811, QN => n1021);
   REGISTERS_reg_29_17_inst : DFFR_X1 port map( D => n7259, CK => CLK, RN => 
                           n3162, Q => n9812, QN => n1022);
   REGISTERS_reg_29_16_inst : DFFR_X1 port map( D => n7260, CK => CLK, RN => 
                           n3162, Q => n9813, QN => n1023);
   REGISTERS_reg_29_15_inst : DFFR_X1 port map( D => n7261, CK => CLK, RN => 
                           n3162, Q => n9814, QN => n1024);
   REGISTERS_reg_29_14_inst : DFFR_X1 port map( D => n7262, CK => CLK, RN => 
                           n3162, Q => n9815, QN => n1025);
   REGISTERS_reg_29_13_inst : DFFR_X1 port map( D => n7263, CK => CLK, RN => 
                           n3162, Q => n9816, QN => n1026);
   REGISTERS_reg_29_12_inst : DFFR_X1 port map( D => n7264, CK => CLK, RN => 
                           n3162, Q => n9817, QN => n1027);
   REGISTERS_reg_29_11_inst : DFFR_X1 port map( D => n7265, CK => CLK, RN => 
                           n3162, Q => n9818, QN => n1028);
   REGISTERS_reg_29_10_inst : DFFR_X1 port map( D => n7266, CK => CLK, RN => 
                           n3162, Q => n9819, QN => n1029);
   REGISTERS_reg_29_9_inst : DFFR_X1 port map( D => n7267, CK => CLK, RN => 
                           n3162, Q => n9820, QN => n1030);
   REGISTERS_reg_29_8_inst : DFFR_X1 port map( D => n7268, CK => CLK, RN => 
                           n3162, Q => n9821, QN => n1031);
   REGISTERS_reg_29_7_inst : DFFR_X1 port map( D => n7269, CK => CLK, RN => 
                           n3160, Q => n9822, QN => n1032);
   REGISTERS_reg_29_6_inst : DFFR_X1 port map( D => n7270, CK => CLK, RN => 
                           n3160, Q => n9823, QN => n1033);
   REGISTERS_reg_29_5_inst : DFFR_X1 port map( D => n7271, CK => CLK, RN => 
                           n3160, Q => n9824, QN => n1034);
   REGISTERS_reg_29_4_inst : DFFR_X1 port map( D => n7272, CK => CLK, RN => 
                           n3160, Q => n9825, QN => n1035);
   REGISTERS_reg_29_3_inst : DFFR_X1 port map( D => n7273, CK => CLK, RN => 
                           n3160, Q => n9826, QN => n1036);
   REGISTERS_reg_29_2_inst : DFFR_X1 port map( D => n7274, CK => CLK, RN => 
                           n3160, Q => n9827, QN => n1037);
   REGISTERS_reg_29_1_inst : DFFR_X1 port map( D => n7275, CK => CLK, RN => 
                           n3160, Q => n9828, QN => n1038);
   REGISTERS_reg_29_0_inst : DFFR_X1 port map( D => n7276, CK => CLK, RN => 
                           n3160, Q => n9829, QN => n1039);
   REGISTERS_reg_30_31_inst : DFFR_X1 port map( D => n7277, CK => CLK, RN => 
                           n3160, Q => n9830, QN => n1040);
   REGISTERS_reg_30_30_inst : DFFR_X1 port map( D => n7278, CK => CLK, RN => 
                           n3160, Q => n9831, QN => n1041);
   REGISTERS_reg_30_29_inst : DFFR_X1 port map( D => n7279, CK => CLK, RN => 
                           n3160, Q => n9832, QN => n1042);
   REGISTERS_reg_30_28_inst : DFFR_X1 port map( D => n7280, CK => CLK, RN => 
                           n3160, Q => n9833, QN => n1043);
   REGISTERS_reg_30_27_inst : DFFR_X1 port map( D => n7281, CK => CLK, RN => 
                           n3159, Q => n9834, QN => n1044);
   REGISTERS_reg_30_26_inst : DFFR_X1 port map( D => n7282, CK => CLK, RN => 
                           n3159, Q => n9835, QN => n1045);
   REGISTERS_reg_30_25_inst : DFFR_X1 port map( D => n7283, CK => CLK, RN => 
                           n3159, Q => n9836, QN => n1046);
   REGISTERS_reg_30_24_inst : DFFR_X1 port map( D => n7284, CK => CLK, RN => 
                           n3159, Q => n9837, QN => n1047);
   REGISTERS_reg_30_23_inst : DFFR_X1 port map( D => n7285, CK => CLK, RN => 
                           n3159, Q => n9838, QN => n1048);
   REGISTERS_reg_30_22_inst : DFFR_X1 port map( D => n7286, CK => CLK, RN => 
                           n3159, Q => n9839, QN => n1049);
   REGISTERS_reg_30_21_inst : DFFR_X1 port map( D => n7287, CK => CLK, RN => 
                           n3159, Q => n9840, QN => n1050);
   REGISTERS_reg_30_20_inst : DFFR_X1 port map( D => n7288, CK => CLK, RN => 
                           n3159, Q => n9841, QN => n1051);
   REGISTERS_reg_30_19_inst : DFFR_X1 port map( D => n7289, CK => CLK, RN => 
                           n3159, Q => n9842, QN => n1052);
   REGISTERS_reg_30_18_inst : DFFR_X1 port map( D => n7290, CK => CLK, RN => 
                           n3159, Q => n9843, QN => n1053);
   REGISTERS_reg_30_17_inst : DFFR_X1 port map( D => n7291, CK => CLK, RN => 
                           n3159, Q => n9844, QN => n1054);
   REGISTERS_reg_30_16_inst : DFFR_X1 port map( D => n7292, CK => CLK, RN => 
                           n3159, Q => n9845, QN => n1055);
   REGISTERS_reg_30_15_inst : DFFR_X1 port map( D => n7293, CK => CLK, RN => 
                           n3158, Q => n9846, QN => n1056);
   REGISTERS_reg_30_14_inst : DFFR_X1 port map( D => n7294, CK => CLK, RN => 
                           n3158, Q => n9847, QN => n1057);
   REGISTERS_reg_30_13_inst : DFFR_X1 port map( D => n7295, CK => CLK, RN => 
                           n3158, Q => n9848, QN => n1058);
   REGISTERS_reg_30_12_inst : DFFR_X1 port map( D => n7296, CK => CLK, RN => 
                           n3158, Q => n9849, QN => n1059);
   REGISTERS_reg_30_11_inst : DFFR_X1 port map( D => n7297, CK => CLK, RN => 
                           n3158, Q => n9850, QN => n1060);
   REGISTERS_reg_30_10_inst : DFFR_X1 port map( D => n7298, CK => CLK, RN => 
                           n3158, Q => n9851, QN => n1061);
   REGISTERS_reg_30_9_inst : DFFR_X1 port map( D => n7299, CK => CLK, RN => 
                           n3158, Q => n9852, QN => n1062);
   REGISTERS_reg_30_8_inst : DFFR_X1 port map( D => n7300, CK => CLK, RN => 
                           n3158, Q => n9853, QN => n1063);
   REGISTERS_reg_30_7_inst : DFFR_X1 port map( D => n7301, CK => CLK, RN => 
                           n3158, Q => n9854, QN => n1064);
   REGISTERS_reg_30_6_inst : DFFR_X1 port map( D => n7302, CK => CLK, RN => 
                           n3158, Q => n9855, QN => n1065);
   REGISTERS_reg_30_5_inst : DFFR_X1 port map( D => n7303, CK => CLK, RN => 
                           n3158, Q => n9856, QN => n1066);
   REGISTERS_reg_30_4_inst : DFFR_X1 port map( D => n7304, CK => CLK, RN => 
                           n3158, Q => n9857, QN => n1067);
   REGISTERS_reg_30_3_inst : DFFR_X1 port map( D => n7305, CK => CLK, RN => 
                           n3156, Q => n9858, QN => n1068);
   REGISTERS_reg_30_2_inst : DFFR_X1 port map( D => n7306, CK => CLK, RN => 
                           n3156, Q => n9859, QN => n1069);
   REGISTERS_reg_30_1_inst : DFFR_X1 port map( D => n7307, CK => CLK, RN => 
                           n3156, Q => n9860, QN => n1070);
   REGISTERS_reg_30_0_inst : DFFR_X1 port map( D => n7308, CK => CLK, RN => 
                           n3156, Q => n9861, QN => n1071);
   REGISTERS_reg_31_31_inst : DFFR_X1 port map( D => n7309, CK => CLK, RN => 
                           n3156, Q => n9862, QN => n1072);
   REGISTERS_reg_31_30_inst : DFFR_X1 port map( D => n7310, CK => CLK, RN => 
                           n3156, Q => n9863, QN => n1073);
   REGISTERS_reg_31_29_inst : DFFR_X1 port map( D => n7311, CK => CLK, RN => 
                           n3156, Q => n9864, QN => n1074);
   REGISTERS_reg_31_28_inst : DFFR_X1 port map( D => n7312, CK => CLK, RN => 
                           n3156, Q => n9865, QN => n1075);
   REGISTERS_reg_31_27_inst : DFFR_X1 port map( D => n7313, CK => CLK, RN => 
                           n3156, Q => n9866, QN => n1076);
   REGISTERS_reg_31_26_inst : DFFR_X1 port map( D => n7314, CK => CLK, RN => 
                           n3156, Q => n9867, QN => n1077);
   REGISTERS_reg_31_25_inst : DFFR_X1 port map( D => n7315, CK => CLK, RN => 
                           n3156, Q => n9868, QN => n1078);
   REGISTERS_reg_31_24_inst : DFFR_X1 port map( D => n7316, CK => CLK, RN => 
                           n3156, Q => n9869, QN => n1079);
   REGISTERS_reg_31_23_inst : DFFR_X1 port map( D => n7317, CK => CLK, RN => 
                           n3155, Q => n9870, QN => n1080);
   REGISTERS_reg_31_22_inst : DFFR_X1 port map( D => n7318, CK => CLK, RN => 
                           n3155, Q => n9871, QN => n1081);
   REGISTERS_reg_31_21_inst : DFFR_X1 port map( D => n7319, CK => CLK, RN => 
                           n3155, Q => n9872, QN => n1082);
   REGISTERS_reg_31_20_inst : DFFR_X1 port map( D => n7320, CK => CLK, RN => 
                           n3155, Q => n9873, QN => n1083);
   REGISTERS_reg_31_19_inst : DFFR_X1 port map( D => n7321, CK => CLK, RN => 
                           n3155, Q => n9874, QN => n1084);
   REGISTERS_reg_31_18_inst : DFFR_X1 port map( D => n7322, CK => CLK, RN => 
                           n3155, Q => n9875, QN => n1085);
   REGISTERS_reg_31_17_inst : DFFR_X1 port map( D => n7323, CK => CLK, RN => 
                           n3155, Q => n9876, QN => n1086);
   REGISTERS_reg_31_16_inst : DFFR_X1 port map( D => n7324, CK => CLK, RN => 
                           n3155, Q => n9877, QN => n1087);
   REGISTERS_reg_31_15_inst : DFFR_X1 port map( D => n7325, CK => CLK, RN => 
                           n3155, Q => n9878, QN => n1088);
   REGISTERS_reg_31_14_inst : DFFR_X1 port map( D => n7326, CK => CLK, RN => 
                           n3155, Q => n9879, QN => n1089);
   REGISTERS_reg_31_13_inst : DFFR_X1 port map( D => n7327, CK => CLK, RN => 
                           n3155, Q => n9880, QN => n1090);
   REGISTERS_reg_31_12_inst : DFFR_X1 port map( D => n7328, CK => CLK, RN => 
                           n3155, Q => n9881, QN => n1091);
   REGISTERS_reg_31_11_inst : DFFR_X1 port map( D => n7329, CK => CLK, RN => 
                           n3154, Q => n9882, QN => n1092);
   REGISTERS_reg_31_10_inst : DFFR_X1 port map( D => n7330, CK => CLK, RN => 
                           n3154, Q => n9883, QN => n1093);
   REGISTERS_reg_31_9_inst : DFFR_X1 port map( D => n7331, CK => CLK, RN => 
                           n3154, Q => n9884, QN => n1094);
   REGISTERS_reg_31_8_inst : DFFR_X1 port map( D => n7332, CK => CLK, RN => 
                           n3154, Q => n9885, QN => n1095);
   REGISTERS_reg_31_7_inst : DFFR_X1 port map( D => n7333, CK => CLK, RN => 
                           n3154, Q => n9886, QN => n1096);
   REGISTERS_reg_31_6_inst : DFFR_X1 port map( D => n7334, CK => CLK, RN => 
                           n3154, Q => n9887, QN => n1097);
   REGISTERS_reg_31_5_inst : DFFR_X1 port map( D => n7335, CK => CLK, RN => 
                           n3154, Q => n9888, QN => n1098);
   REGISTERS_reg_31_4_inst : DFFR_X1 port map( D => n7336, CK => CLK, RN => 
                           n3154, Q => n9889, QN => n1099);
   REGISTERS_reg_31_3_inst : DFFR_X1 port map( D => n7337, CK => CLK, RN => 
                           n3154, Q => n9890, QN => n1100);
   REGISTERS_reg_31_2_inst : DFFR_X1 port map( D => n7338, CK => CLK, RN => 
                           n3154, Q => n9891, QN => n1101);
   REGISTERS_reg_31_1_inst : DFFR_X1 port map( D => n7339, CK => CLK, RN => 
                           n3154, Q => n9892, QN => n1102);
   REGISTERS_reg_31_0_inst : DFFR_X1 port map( D => n7340, CK => CLK, RN => 
                           n3154, Q => n9893, QN => n1103);
   REGISTERS_reg_32_31_inst : DFFR_X1 port map( D => n7341, CK => CLK, RN => 
                           n3152, Q => n9894, QN => n1104);
   REGISTERS_reg_32_30_inst : DFFR_X1 port map( D => n7342, CK => CLK, RN => 
                           n3152, Q => n9895, QN => n1105);
   REGISTERS_reg_32_29_inst : DFFR_X1 port map( D => n7343, CK => CLK, RN => 
                           n3152, Q => n9896, QN => n1106);
   REGISTERS_reg_32_28_inst : DFFR_X1 port map( D => n7344, CK => CLK, RN => 
                           n3152, Q => n9897, QN => n1107);
   REGISTERS_reg_32_27_inst : DFFR_X1 port map( D => n7345, CK => CLK, RN => 
                           n3152, Q => n9898, QN => n1108);
   REGISTERS_reg_32_26_inst : DFFR_X1 port map( D => n7346, CK => CLK, RN => 
                           n3152, Q => n9899, QN => n1109);
   REGISTERS_reg_32_25_inst : DFFR_X1 port map( D => n7347, CK => CLK, RN => 
                           n3152, Q => n9900, QN => n1110);
   REGISTERS_reg_32_24_inst : DFFR_X1 port map( D => n7348, CK => CLK, RN => 
                           n3152, Q => n9901, QN => n1111);
   REGISTERS_reg_32_23_inst : DFFR_X1 port map( D => n7349, CK => CLK, RN => 
                           n3152, Q => n9902, QN => n1112);
   REGISTERS_reg_32_22_inst : DFFR_X1 port map( D => n7350, CK => CLK, RN => 
                           n3152, Q => n9903, QN => n1113);
   REGISTERS_reg_32_21_inst : DFFR_X1 port map( D => n7351, CK => CLK, RN => 
                           n3152, Q => n9904, QN => n1114);
   REGISTERS_reg_32_20_inst : DFFR_X1 port map( D => n7352, CK => CLK, RN => 
                           n3152, Q => n9905, QN => n1115);
   REGISTERS_reg_32_19_inst : DFFR_X1 port map( D => n7353, CK => CLK, RN => 
                           n3151, Q => n9906, QN => n1116);
   REGISTERS_reg_32_18_inst : DFFR_X1 port map( D => n7354, CK => CLK, RN => 
                           n3151, Q => n9907, QN => n1117);
   REGISTERS_reg_32_17_inst : DFFR_X1 port map( D => n7355, CK => CLK, RN => 
                           n3151, Q => n9908, QN => n1118);
   REGISTERS_reg_32_16_inst : DFFR_X1 port map( D => n7356, CK => CLK, RN => 
                           n3151, Q => n9909, QN => n1119);
   REGISTERS_reg_32_15_inst : DFFR_X1 port map( D => n7357, CK => CLK, RN => 
                           n3151, Q => n9910, QN => n1120);
   REGISTERS_reg_32_14_inst : DFFR_X1 port map( D => n7358, CK => CLK, RN => 
                           n3151, Q => n9911, QN => n1121);
   REGISTERS_reg_32_13_inst : DFFR_X1 port map( D => n7359, CK => CLK, RN => 
                           n3151, Q => n9912, QN => n1122);
   REGISTERS_reg_32_12_inst : DFFR_X1 port map( D => n7360, CK => CLK, RN => 
                           n3151, Q => n9913, QN => n1123);
   REGISTERS_reg_32_11_inst : DFFR_X1 port map( D => n7361, CK => CLK, RN => 
                           n3151, Q => n9914, QN => n1124);
   REGISTERS_reg_32_10_inst : DFFR_X1 port map( D => n7362, CK => CLK, RN => 
                           n3151, Q => n9915, QN => n1125);
   REGISTERS_reg_32_9_inst : DFFR_X1 port map( D => n7363, CK => CLK, RN => 
                           n3151, Q => n9916, QN => n1126);
   REGISTERS_reg_32_8_inst : DFFR_X1 port map( D => n7364, CK => CLK, RN => 
                           n3151, Q => n9917, QN => n1127);
   REGISTERS_reg_32_7_inst : DFFR_X1 port map( D => n7365, CK => CLK, RN => 
                           n3150, Q => n9918, QN => n1128);
   REGISTERS_reg_32_6_inst : DFFR_X1 port map( D => n7366, CK => CLK, RN => 
                           n3150, Q => n9919, QN => n1129);
   REGISTERS_reg_32_5_inst : DFFR_X1 port map( D => n7367, CK => CLK, RN => 
                           n3150, Q => n9920, QN => n1130);
   REGISTERS_reg_32_4_inst : DFFR_X1 port map( D => n7368, CK => CLK, RN => 
                           n3150, Q => n9921, QN => n1131);
   REGISTERS_reg_32_3_inst : DFFR_X1 port map( D => n7369, CK => CLK, RN => 
                           n3150, Q => n9922, QN => n1132);
   REGISTERS_reg_32_2_inst : DFFR_X1 port map( D => n7370, CK => CLK, RN => 
                           n3150, Q => n9923, QN => n1133);
   REGISTERS_reg_32_1_inst : DFFR_X1 port map( D => n7371, CK => CLK, RN => 
                           n3150, Q => n9924, QN => n1134);
   REGISTERS_reg_32_0_inst : DFFR_X1 port map( D => n7372, CK => CLK, RN => 
                           n3150, Q => n9925, QN => n1135);
   REGISTERS_reg_35_31_inst : DFFR_X1 port map( D => n7437, CK => CLK, RN => 
                           n3142, Q => n9926, QN => n1200);
   REGISTERS_reg_35_30_inst : DFFR_X1 port map( D => n7438, CK => CLK, RN => 
                           n3142, Q => n9927, QN => n1201);
   REGISTERS_reg_35_29_inst : DFFR_X1 port map( D => n7439, CK => CLK, RN => 
                           n3142, Q => n9928, QN => n1202);
   REGISTERS_reg_35_28_inst : DFFR_X1 port map( D => n7440, CK => CLK, RN => 
                           n3142, Q => n9929, QN => n1203);
   REGISTERS_reg_35_27_inst : DFFR_X1 port map( D => n7441, CK => CLK, RN => 
                           n3142, Q => n9930, QN => n1204);
   REGISTERS_reg_35_26_inst : DFFR_X1 port map( D => n7442, CK => CLK, RN => 
                           n3142, Q => n9931, QN => n1205);
   REGISTERS_reg_35_25_inst : DFFR_X1 port map( D => n7443, CK => CLK, RN => 
                           n3142, Q => n9932, QN => n1206);
   REGISTERS_reg_35_24_inst : DFFR_X1 port map( D => n7444, CK => CLK, RN => 
                           n3142, Q => n9933, QN => n1207);
   REGISTERS_reg_35_23_inst : DFFR_X1 port map( D => n7445, CK => CLK, RN => 
                           n3142, Q => n9934, QN => n1208);
   REGISTERS_reg_35_22_inst : DFFR_X1 port map( D => n7446, CK => CLK, RN => 
                           n3142, Q => n9935, QN => n1209);
   REGISTERS_reg_35_21_inst : DFFR_X1 port map( D => n7447, CK => CLK, RN => 
                           n3142, Q => n9936, QN => n1210);
   REGISTERS_reg_35_20_inst : DFFR_X1 port map( D => n7448, CK => CLK, RN => 
                           n3142, Q => n9937, QN => n1211);
   REGISTERS_reg_35_19_inst : DFFR_X1 port map( D => n7449, CK => CLK, RN => 
                           n3140, Q => n9938, QN => n1212);
   REGISTERS_reg_35_18_inst : DFFR_X1 port map( D => n7450, CK => CLK, RN => 
                           n3140, Q => n9939, QN => n1213);
   REGISTERS_reg_35_17_inst : DFFR_X1 port map( D => n7451, CK => CLK, RN => 
                           n3140, Q => n9940, QN => n1214);
   REGISTERS_reg_35_16_inst : DFFR_X1 port map( D => n7452, CK => CLK, RN => 
                           n3140, Q => n9941, QN => n1215);
   REGISTERS_reg_35_15_inst : DFFR_X1 port map( D => n7453, CK => CLK, RN => 
                           n3140, Q => n9942, QN => n1216);
   REGISTERS_reg_35_14_inst : DFFR_X1 port map( D => n7454, CK => CLK, RN => 
                           n3140, Q => n9943, QN => n1217);
   REGISTERS_reg_35_13_inst : DFFR_X1 port map( D => n7455, CK => CLK, RN => 
                           n3140, Q => n9944, QN => n1218);
   REGISTERS_reg_35_12_inst : DFFR_X1 port map( D => n7456, CK => CLK, RN => 
                           n3140, Q => n9945, QN => n1219);
   REGISTERS_reg_35_11_inst : DFFR_X1 port map( D => n7457, CK => CLK, RN => 
                           n3140, Q => n9946, QN => n1220);
   REGISTERS_reg_35_10_inst : DFFR_X1 port map( D => n7458, CK => CLK, RN => 
                           n3140, Q => n9947, QN => n1221);
   REGISTERS_reg_35_9_inst : DFFR_X1 port map( D => n7459, CK => CLK, RN => 
                           n3140, Q => n9948, QN => n1222);
   REGISTERS_reg_35_8_inst : DFFR_X1 port map( D => n7460, CK => CLK, RN => 
                           n3140, Q => n9949, QN => n1223);
   REGISTERS_reg_35_7_inst : DFFR_X1 port map( D => n7461, CK => CLK, RN => 
                           n3139, Q => n9950, QN => n1224);
   REGISTERS_reg_35_6_inst : DFFR_X1 port map( D => n7462, CK => CLK, RN => 
                           n3139, Q => n9951, QN => n1225);
   REGISTERS_reg_35_5_inst : DFFR_X1 port map( D => n7463, CK => CLK, RN => 
                           n3139, Q => n9952, QN => n1226);
   REGISTERS_reg_35_4_inst : DFFR_X1 port map( D => n7464, CK => CLK, RN => 
                           n3139, Q => n9953, QN => n1227);
   REGISTERS_reg_35_3_inst : DFFR_X1 port map( D => n7465, CK => CLK, RN => 
                           n3139, Q => n9954, QN => n1228);
   REGISTERS_reg_35_2_inst : DFFR_X1 port map( D => n7466, CK => CLK, RN => 
                           n3139, Q => n9955, QN => n1229);
   REGISTERS_reg_35_1_inst : DFFR_X1 port map( D => n7467, CK => CLK, RN => 
                           n3139, Q => n9956, QN => n1230);
   REGISTERS_reg_35_0_inst : DFFR_X1 port map( D => n7468, CK => CLK, RN => 
                           n3139, Q => n9957, QN => n1231);
   REGISTERS_reg_36_31_inst : DFFR_X1 port map( D => n7469, CK => CLK, RN => 
                           n3139, Q => n9958, QN => n1232);
   REGISTERS_reg_36_30_inst : DFFR_X1 port map( D => n7470, CK => CLK, RN => 
                           n3139, Q => n9959, QN => n1233);
   REGISTERS_reg_36_29_inst : DFFR_X1 port map( D => n7471, CK => CLK, RN => 
                           n3139, Q => n9960, QN => n1234);
   REGISTERS_reg_36_28_inst : DFFR_X1 port map( D => n7472, CK => CLK, RN => 
                           n3139, Q => n9961, QN => n1235);
   REGISTERS_reg_36_27_inst : DFFR_X1 port map( D => n7473, CK => CLK, RN => 
                           n3138, Q => n9962, QN => n1236);
   REGISTERS_reg_36_26_inst : DFFR_X1 port map( D => n7474, CK => CLK, RN => 
                           n3138, Q => n9963, QN => n1237);
   REGISTERS_reg_36_25_inst : DFFR_X1 port map( D => n7475, CK => CLK, RN => 
                           n3138, Q => n9964, QN => n1238);
   REGISTERS_reg_36_24_inst : DFFR_X1 port map( D => n7476, CK => CLK, RN => 
                           n3138, Q => n9965, QN => n1239);
   REGISTERS_reg_36_23_inst : DFFR_X1 port map( D => n7477, CK => CLK, RN => 
                           n3138, Q => n9966, QN => n1240);
   REGISTERS_reg_36_22_inst : DFFR_X1 port map( D => n7478, CK => CLK, RN => 
                           n3138, Q => n9967, QN => n1241);
   REGISTERS_reg_36_21_inst : DFFR_X1 port map( D => n7479, CK => CLK, RN => 
                           n3138, Q => n9968, QN => n1242);
   REGISTERS_reg_36_20_inst : DFFR_X1 port map( D => n7480, CK => CLK, RN => 
                           n3138, Q => n9969, QN => n1243);
   REGISTERS_reg_36_19_inst : DFFR_X1 port map( D => n7481, CK => CLK, RN => 
                           n3138, Q => n9970, QN => n1244);
   REGISTERS_reg_36_18_inst : DFFR_X1 port map( D => n7482, CK => CLK, RN => 
                           n3138, Q => n9971, QN => n1245);
   REGISTERS_reg_36_17_inst : DFFR_X1 port map( D => n7483, CK => CLK, RN => 
                           n3138, Q => n9972, QN => n1246);
   REGISTERS_reg_36_16_inst : DFFR_X1 port map( D => n7484, CK => CLK, RN => 
                           n3138, Q => n9973, QN => n1247);
   REGISTERS_reg_36_15_inst : DFFR_X1 port map( D => n7485, CK => CLK, RN => 
                           n3136, Q => n9974, QN => n1248);
   REGISTERS_reg_36_14_inst : DFFR_X1 port map( D => n7486, CK => CLK, RN => 
                           n3136, Q => n9975, QN => n1249);
   REGISTERS_reg_36_13_inst : DFFR_X1 port map( D => n7487, CK => CLK, RN => 
                           n3136, Q => n9976, QN => n1250);
   REGISTERS_reg_36_12_inst : DFFR_X1 port map( D => n7488, CK => CLK, RN => 
                           n3136, Q => n9977, QN => n1251);
   REGISTERS_reg_36_11_inst : DFFR_X1 port map( D => n7489, CK => CLK, RN => 
                           n3136, Q => n9978, QN => n1252);
   REGISTERS_reg_36_10_inst : DFFR_X1 port map( D => n7490, CK => CLK, RN => 
                           n3136, Q => n9979, QN => n1253);
   REGISTERS_reg_36_9_inst : DFFR_X1 port map( D => n7491, CK => CLK, RN => 
                           n3136, Q => n9980, QN => n1254);
   REGISTERS_reg_36_8_inst : DFFR_X1 port map( D => n7492, CK => CLK, RN => 
                           n3136, Q => n9981, QN => n1255);
   REGISTERS_reg_36_7_inst : DFFR_X1 port map( D => n7493, CK => CLK, RN => 
                           n3136, Q => n9982, QN => n1256);
   REGISTERS_reg_36_6_inst : DFFR_X1 port map( D => n7494, CK => CLK, RN => 
                           n3136, Q => n9983, QN => n1257);
   REGISTERS_reg_36_5_inst : DFFR_X1 port map( D => n7495, CK => CLK, RN => 
                           n3136, Q => n9984, QN => n1258);
   REGISTERS_reg_36_4_inst : DFFR_X1 port map( D => n7496, CK => CLK, RN => 
                           n3136, Q => n9985, QN => n1259);
   REGISTERS_reg_36_3_inst : DFFR_X1 port map( D => n7497, CK => CLK, RN => 
                           n3135, Q => n9986, QN => n1260);
   REGISTERS_reg_36_2_inst : DFFR_X1 port map( D => n7498, CK => CLK, RN => 
                           n3135, Q => n9987, QN => n1261);
   REGISTERS_reg_36_1_inst : DFFR_X1 port map( D => n7499, CK => CLK, RN => 
                           n3135, Q => n9988, QN => n1262);
   REGISTERS_reg_36_0_inst : DFFR_X1 port map( D => n7500, CK => CLK, RN => 
                           n3135, Q => n9989, QN => n1263);
   REGISTERS_reg_37_31_inst : DFFR_X1 port map( D => n7501, CK => CLK, RN => 
                           n3135, Q => n9990, QN => n1264);
   REGISTERS_reg_37_30_inst : DFFR_X1 port map( D => n7502, CK => CLK, RN => 
                           n3135, Q => n9991, QN => n1265);
   REGISTERS_reg_37_29_inst : DFFR_X1 port map( D => n7503, CK => CLK, RN => 
                           n3135, Q => n9992, QN => n1266);
   REGISTERS_reg_37_28_inst : DFFR_X1 port map( D => n7504, CK => CLK, RN => 
                           n3135, Q => n9993, QN => n1267);
   REGISTERS_reg_37_27_inst : DFFR_X1 port map( D => n7505, CK => CLK, RN => 
                           n3135, Q => n9994, QN => n1268);
   REGISTERS_reg_37_26_inst : DFFR_X1 port map( D => n7506, CK => CLK, RN => 
                           n3135, Q => n9995, QN => n1269);
   REGISTERS_reg_37_25_inst : DFFR_X1 port map( D => n7507, CK => CLK, RN => 
                           n3135, Q => n9996, QN => n1270);
   REGISTERS_reg_37_24_inst : DFFR_X1 port map( D => n7508, CK => CLK, RN => 
                           n3135, Q => n9997, QN => n1271);
   REGISTERS_reg_37_23_inst : DFFR_X1 port map( D => n7509, CK => CLK, RN => 
                           n3134, Q => n9998, QN => n1272);
   REGISTERS_reg_37_22_inst : DFFR_X1 port map( D => n7510, CK => CLK, RN => 
                           n3134, Q => n9999, QN => n1273);
   REGISTERS_reg_37_21_inst : DFFR_X1 port map( D => n7511, CK => CLK, RN => 
                           n3134, Q => n10000, QN => n1274);
   REGISTERS_reg_37_20_inst : DFFR_X1 port map( D => n7512, CK => CLK, RN => 
                           n3134, Q => n10001, QN => n1275);
   REGISTERS_reg_37_19_inst : DFFR_X1 port map( D => n7513, CK => CLK, RN => 
                           n3134, Q => n10002, QN => n1276);
   REGISTERS_reg_37_18_inst : DFFR_X1 port map( D => n7514, CK => CLK, RN => 
                           n3134, Q => n10003, QN => n1277);
   REGISTERS_reg_37_17_inst : DFFR_X1 port map( D => n7515, CK => CLK, RN => 
                           n3134, Q => n10004, QN => n1278);
   REGISTERS_reg_37_16_inst : DFFR_X1 port map( D => n7516, CK => CLK, RN => 
                           n3134, Q => n10005, QN => n1279);
   REGISTERS_reg_37_15_inst : DFFR_X1 port map( D => n7517, CK => CLK, RN => 
                           n3134, Q => n10006, QN => n1280);
   REGISTERS_reg_37_14_inst : DFFR_X1 port map( D => n7518, CK => CLK, RN => 
                           n3134, Q => n10007, QN => n1281);
   REGISTERS_reg_37_13_inst : DFFR_X1 port map( D => n7519, CK => CLK, RN => 
                           n3134, Q => n10008, QN => n1282);
   REGISTERS_reg_37_12_inst : DFFR_X1 port map( D => n7520, CK => CLK, RN => 
                           n3134, Q => n10009, QN => n1283);
   REGISTERS_reg_37_11_inst : DFFR_X1 port map( D => n7521, CK => CLK, RN => 
                           n3132, Q => n10010, QN => n1284);
   REGISTERS_reg_37_10_inst : DFFR_X1 port map( D => n7522, CK => CLK, RN => 
                           n3132, Q => n10011, QN => n1285);
   REGISTERS_reg_37_9_inst : DFFR_X1 port map( D => n7523, CK => CLK, RN => 
                           n3132, Q => n10012, QN => n1286);
   REGISTERS_reg_37_8_inst : DFFR_X1 port map( D => n7524, CK => CLK, RN => 
                           n3132, Q => n10013, QN => n1287);
   REGISTERS_reg_37_7_inst : DFFR_X1 port map( D => n7525, CK => CLK, RN => 
                           n3132, Q => n10014, QN => n1288);
   REGISTERS_reg_37_6_inst : DFFR_X1 port map( D => n7526, CK => CLK, RN => 
                           n3132, Q => n10015, QN => n1289);
   REGISTERS_reg_37_5_inst : DFFR_X1 port map( D => n7527, CK => CLK, RN => 
                           n3132, Q => n10016, QN => n1290);
   REGISTERS_reg_37_4_inst : DFFR_X1 port map( D => n7528, CK => CLK, RN => 
                           n3132, Q => n10017, QN => n1291);
   REGISTERS_reg_37_3_inst : DFFR_X1 port map( D => n7529, CK => CLK, RN => 
                           n3132, Q => n10018, QN => n1292);
   REGISTERS_reg_37_2_inst : DFFR_X1 port map( D => n7530, CK => CLK, RN => 
                           n3132, Q => n10019, QN => n1293);
   REGISTERS_reg_37_1_inst : DFFR_X1 port map( D => n7531, CK => CLK, RN => 
                           n3132, Q => n10020, QN => n1294);
   REGISTERS_reg_37_0_inst : DFFR_X1 port map( D => n7532, CK => CLK, RN => 
                           n3132, Q => n10021, QN => n1295);
   REGISTERS_reg_46_31_inst : DFFR_X1 port map( D => n7789, CK => CLK, RN => 
                           n3096, Q => n10022, QN => n1552);
   REGISTERS_reg_46_30_inst : DFFR_X1 port map( D => n7790, CK => CLK, RN => 
                           n3096, Q => n10023, QN => n1553);
   REGISTERS_reg_46_29_inst : DFFR_X1 port map( D => n7791, CK => CLK, RN => 
                           n3096, Q => n10024, QN => n1554);
   REGISTERS_reg_46_28_inst : DFFR_X1 port map( D => n7792, CK => CLK, RN => 
                           n3096, Q => n10025, QN => n1555);
   REGISTERS_reg_46_27_inst : DFFR_X1 port map( D => n7793, CK => CLK, RN => 
                           n3096, Q => n10026, QN => n1556);
   REGISTERS_reg_46_26_inst : DFFR_X1 port map( D => n7794, CK => CLK, RN => 
                           n3096, Q => n10027, QN => n1557);
   REGISTERS_reg_46_25_inst : DFFR_X1 port map( D => n7795, CK => CLK, RN => 
                           n3096, Q => n10028, QN => n1558);
   REGISTERS_reg_46_24_inst : DFFR_X1 port map( D => n7796, CK => CLK, RN => 
                           n3096, Q => n10029, QN => n1559);
   REGISTERS_reg_46_23_inst : DFFR_X1 port map( D => n7797, CK => CLK, RN => 
                           n3094, Q => n10030, QN => n1560);
   REGISTERS_reg_46_22_inst : DFFR_X1 port map( D => n7798, CK => CLK, RN => 
                           n3094, Q => n10031, QN => n1561);
   REGISTERS_reg_46_21_inst : DFFR_X1 port map( D => n7799, CK => CLK, RN => 
                           n3094, Q => n10032, QN => n1562);
   REGISTERS_reg_46_20_inst : DFFR_X1 port map( D => n7800, CK => CLK, RN => 
                           n3094, Q => n10033, QN => n1563);
   REGISTERS_reg_46_19_inst : DFFR_X1 port map( D => n7801, CK => CLK, RN => 
                           n3094, Q => n10034, QN => n1564);
   REGISTERS_reg_46_18_inst : DFFR_X1 port map( D => n7802, CK => CLK, RN => 
                           n3094, Q => n10035, QN => n1565);
   REGISTERS_reg_46_17_inst : DFFR_X1 port map( D => n7803, CK => CLK, RN => 
                           n3094, Q => n10036, QN => n1566);
   REGISTERS_reg_46_16_inst : DFFR_X1 port map( D => n7804, CK => CLK, RN => 
                           n3094, Q => n10037, QN => n1567);
   REGISTERS_reg_46_15_inst : DFFR_X1 port map( D => n7805, CK => CLK, RN => 
                           n3094, Q => n10038, QN => n1568);
   REGISTERS_reg_46_14_inst : DFFR_X1 port map( D => n7806, CK => CLK, RN => 
                           n3094, Q => n10039, QN => n1569);
   REGISTERS_reg_46_13_inst : DFFR_X1 port map( D => n7807, CK => CLK, RN => 
                           n3094, Q => n10040, QN => n1570);
   REGISTERS_reg_46_12_inst : DFFR_X1 port map( D => n7808, CK => CLK, RN => 
                           n3094, Q => n10041, QN => n1571);
   REGISTERS_reg_46_11_inst : DFFR_X1 port map( D => n7809, CK => CLK, RN => 
                           n3092, Q => n10042, QN => n1572);
   REGISTERS_reg_46_10_inst : DFFR_X1 port map( D => n7810, CK => CLK, RN => 
                           n3092, Q => n10043, QN => n1573);
   REGISTERS_reg_46_9_inst : DFFR_X1 port map( D => n7811, CK => CLK, RN => 
                           n3092, Q => n10044, QN => n1574);
   REGISTERS_reg_46_8_inst : DFFR_X1 port map( D => n7812, CK => CLK, RN => 
                           n3092, Q => n10045, QN => n1575);
   REGISTERS_reg_46_7_inst : DFFR_X1 port map( D => n7813, CK => CLK, RN => 
                           n3092, Q => n10046, QN => n1576);
   REGISTERS_reg_46_6_inst : DFFR_X1 port map( D => n7814, CK => CLK, RN => 
                           n3092, Q => n10047, QN => n1577);
   REGISTERS_reg_46_5_inst : DFFR_X1 port map( D => n7815, CK => CLK, RN => 
                           n3092, Q => n10048, QN => n1578);
   REGISTERS_reg_46_4_inst : DFFR_X1 port map( D => n7816, CK => CLK, RN => 
                           n3092, Q => n10049, QN => n1579);
   REGISTERS_reg_46_3_inst : DFFR_X1 port map( D => n7817, CK => CLK, RN => 
                           n3092, Q => n10050, QN => n1580);
   REGISTERS_reg_46_2_inst : DFFR_X1 port map( D => n7818, CK => CLK, RN => 
                           n3092, Q => n10051, QN => n1581);
   REGISTERS_reg_46_1_inst : DFFR_X1 port map( D => n7819, CK => CLK, RN => 
                           n3092, Q => n10052, QN => n1582);
   REGISTERS_reg_46_0_inst : DFFR_X1 port map( D => n7820, CK => CLK, RN => 
                           n3092, Q => n10053, QN => n1583);
   REGISTERS_reg_47_31_inst : DFFR_X1 port map( D => n7821, CK => CLK, RN => 
                           n3091, Q => n10054, QN => n1584);
   REGISTERS_reg_47_30_inst : DFFR_X1 port map( D => n7822, CK => CLK, RN => 
                           n3091, Q => n10055, QN => n1585);
   REGISTERS_reg_47_29_inst : DFFR_X1 port map( D => n7823, CK => CLK, RN => 
                           n3091, Q => n10056, QN => n1586);
   REGISTERS_reg_47_28_inst : DFFR_X1 port map( D => n7824, CK => CLK, RN => 
                           n3091, Q => n10057, QN => n1587);
   REGISTERS_reg_47_27_inst : DFFR_X1 port map( D => n7825, CK => CLK, RN => 
                           n3091, Q => n10058, QN => n1588);
   REGISTERS_reg_47_26_inst : DFFR_X1 port map( D => n7826, CK => CLK, RN => 
                           n3091, Q => n10059, QN => n1589);
   REGISTERS_reg_47_25_inst : DFFR_X1 port map( D => n7827, CK => CLK, RN => 
                           n3091, Q => n10060, QN => n1590);
   REGISTERS_reg_47_24_inst : DFFR_X1 port map( D => n7828, CK => CLK, RN => 
                           n3091, Q => n10061, QN => n1591);
   REGISTERS_reg_47_23_inst : DFFR_X1 port map( D => n7829, CK => CLK, RN => 
                           n3091, Q => n10062, QN => n1592);
   REGISTERS_reg_47_22_inst : DFFR_X1 port map( D => n7830, CK => CLK, RN => 
                           n3091, Q => n10063, QN => n1593);
   REGISTERS_reg_47_21_inst : DFFR_X1 port map( D => n7831, CK => CLK, RN => 
                           n3091, Q => n10064, QN => n1594);
   REGISTERS_reg_47_20_inst : DFFR_X1 port map( D => n7832, CK => CLK, RN => 
                           n3091, Q => n10065, QN => n1595);
   REGISTERS_reg_47_19_inst : DFFR_X1 port map( D => n7833, CK => CLK, RN => 
                           n3089, Q => n10066, QN => n1596);
   REGISTERS_reg_47_18_inst : DFFR_X1 port map( D => n7834, CK => CLK, RN => 
                           n3089, Q => n10067, QN => n1597);
   REGISTERS_reg_47_17_inst : DFFR_X1 port map( D => n7835, CK => CLK, RN => 
                           n3089, Q => n10068, QN => n1598);
   REGISTERS_reg_47_16_inst : DFFR_X1 port map( D => n7836, CK => CLK, RN => 
                           n3089, Q => n10069, QN => n1599);
   REGISTERS_reg_47_15_inst : DFFR_X1 port map( D => n7837, CK => CLK, RN => 
                           n3089, Q => n10070, QN => n1600);
   REGISTERS_reg_47_14_inst : DFFR_X1 port map( D => n7838, CK => CLK, RN => 
                           n3089, Q => n10071, QN => n1601);
   REGISTERS_reg_47_13_inst : DFFR_X1 port map( D => n7839, CK => CLK, RN => 
                           n3089, Q => n10072, QN => n1602);
   REGISTERS_reg_47_12_inst : DFFR_X1 port map( D => n7840, CK => CLK, RN => 
                           n3089, Q => n10073, QN => n1603);
   REGISTERS_reg_47_11_inst : DFFR_X1 port map( D => n7841, CK => CLK, RN => 
                           n3089, Q => n10074, QN => n1604);
   REGISTERS_reg_47_10_inst : DFFR_X1 port map( D => n7842, CK => CLK, RN => 
                           n3089, Q => n10075, QN => n1605);
   REGISTERS_reg_47_9_inst : DFFR_X1 port map( D => n7843, CK => CLK, RN => 
                           n3089, Q => n10076, QN => n1606);
   REGISTERS_reg_47_8_inst : DFFR_X1 port map( D => n7844, CK => CLK, RN => 
                           n3089, Q => n10077, QN => n1607);
   REGISTERS_reg_47_7_inst : DFFR_X1 port map( D => n7845, CK => CLK, RN => 
                           n3087, Q => n10078, QN => n1608);
   REGISTERS_reg_47_6_inst : DFFR_X1 port map( D => n7846, CK => CLK, RN => 
                           n3087, Q => n10079, QN => n1609);
   REGISTERS_reg_47_5_inst : DFFR_X1 port map( D => n7847, CK => CLK, RN => 
                           n3087, Q => n10080, QN => n1610);
   REGISTERS_reg_47_4_inst : DFFR_X1 port map( D => n7848, CK => CLK, RN => 
                           n3087, Q => n10081, QN => n1611);
   REGISTERS_reg_47_3_inst : DFFR_X1 port map( D => n7849, CK => CLK, RN => 
                           n3087, Q => n10082, QN => n1612);
   REGISTERS_reg_47_2_inst : DFFR_X1 port map( D => n7850, CK => CLK, RN => 
                           n3087, Q => n10083, QN => n1613);
   REGISTERS_reg_47_1_inst : DFFR_X1 port map( D => n7851, CK => CLK, RN => 
                           n3087, Q => n10084, QN => n1614);
   REGISTERS_reg_47_0_inst : DFFR_X1 port map( D => n7852, CK => CLK, RN => 
                           n3087, Q => n10085, QN => n1615);
   REGISTERS_reg_48_31_inst : DFFR_X1 port map( D => n7853, CK => CLK, RN => 
                           n3087, Q => n10086, QN => n1616);
   REGISTERS_reg_48_30_inst : DFFR_X1 port map( D => n7854, CK => CLK, RN => 
                           n3087, Q => n10087, QN => n1617);
   REGISTERS_reg_48_29_inst : DFFR_X1 port map( D => n7855, CK => CLK, RN => 
                           n3087, Q => n10088, QN => n1618);
   REGISTERS_reg_48_28_inst : DFFR_X1 port map( D => n7856, CK => CLK, RN => 
                           n3087, Q => n10089, QN => n1619);
   REGISTERS_reg_48_27_inst : DFFR_X1 port map( D => n7857, CK => CLK, RN => 
                           n3086, Q => n10090, QN => n1620);
   REGISTERS_reg_48_26_inst : DFFR_X1 port map( D => n7858, CK => CLK, RN => 
                           n3086, Q => n10091, QN => n1621);
   REGISTERS_reg_48_25_inst : DFFR_X1 port map( D => n7859, CK => CLK, RN => 
                           n3086, Q => n10092, QN => n1622);
   REGISTERS_reg_48_24_inst : DFFR_X1 port map( D => n7860, CK => CLK, RN => 
                           n3086, Q => n10093, QN => n1623);
   REGISTERS_reg_48_23_inst : DFFR_X1 port map( D => n7861, CK => CLK, RN => 
                           n3086, Q => n10094, QN => n1624);
   REGISTERS_reg_48_22_inst : DFFR_X1 port map( D => n7862, CK => CLK, RN => 
                           n3086, Q => n10095, QN => n1625);
   REGISTERS_reg_48_21_inst : DFFR_X1 port map( D => n7863, CK => CLK, RN => 
                           n3086, Q => n10096, QN => n1626);
   REGISTERS_reg_48_20_inst : DFFR_X1 port map( D => n7864, CK => CLK, RN => 
                           n3086, Q => n10097, QN => n1627);
   REGISTERS_reg_48_19_inst : DFFR_X1 port map( D => n7865, CK => CLK, RN => 
                           n3086, Q => n10098, QN => n1628);
   REGISTERS_reg_48_18_inst : DFFR_X1 port map( D => n7866, CK => CLK, RN => 
                           n3086, Q => n10099, QN => n1629);
   REGISTERS_reg_48_17_inst : DFFR_X1 port map( D => n7867, CK => CLK, RN => 
                           n3086, Q => n10100, QN => n1630);
   REGISTERS_reg_48_16_inst : DFFR_X1 port map( D => n7868, CK => CLK, RN => 
                           n3086, Q => n10101, QN => n1631);
   REGISTERS_reg_48_15_inst : DFFR_X1 port map( D => n7869, CK => CLK, RN => 
                           n3084, Q => n10102, QN => n1632);
   REGISTERS_reg_48_14_inst : DFFR_X1 port map( D => n7870, CK => CLK, RN => 
                           n3084, Q => n10103, QN => n1633);
   REGISTERS_reg_48_13_inst : DFFR_X1 port map( D => n7871, CK => CLK, RN => 
                           n3084, Q => n10104, QN => n1634);
   REGISTERS_reg_48_12_inst : DFFR_X1 port map( D => n7872, CK => CLK, RN => 
                           n3084, Q => n10105, QN => n1635);
   REGISTERS_reg_48_11_inst : DFFR_X1 port map( D => n7873, CK => CLK, RN => 
                           n3084, Q => n10106, QN => n1636);
   REGISTERS_reg_48_10_inst : DFFR_X1 port map( D => n7874, CK => CLK, RN => 
                           n3084, Q => n10107, QN => n1637);
   REGISTERS_reg_48_9_inst : DFFR_X1 port map( D => n7875, CK => CLK, RN => 
                           n3084, Q => n10108, QN => n1638);
   REGISTERS_reg_48_8_inst : DFFR_X1 port map( D => n7876, CK => CLK, RN => 
                           n3084, Q => n10109, QN => n1639);
   REGISTERS_reg_48_7_inst : DFFR_X1 port map( D => n7877, CK => CLK, RN => 
                           n3084, Q => n10110, QN => n1640);
   REGISTERS_reg_48_6_inst : DFFR_X1 port map( D => n7878, CK => CLK, RN => 
                           n3084, Q => n10111, QN => n1641);
   REGISTERS_reg_48_5_inst : DFFR_X1 port map( D => n7879, CK => CLK, RN => 
                           n3084, Q => n10112, QN => n1642);
   REGISTERS_reg_48_4_inst : DFFR_X1 port map( D => n7880, CK => CLK, RN => 
                           n3084, Q => n10113, QN => n1643);
   REGISTERS_reg_48_3_inst : DFFR_X1 port map( D => n7881, CK => CLK, RN => 
                           n3082, Q => n10114, QN => n1644);
   REGISTERS_reg_48_2_inst : DFFR_X1 port map( D => n7882, CK => CLK, RN => 
                           n3082, Q => n10115, QN => n1645);
   REGISTERS_reg_48_1_inst : DFFR_X1 port map( D => n7883, CK => CLK, RN => 
                           n3082, Q => n10116, QN => n1646);
   REGISTERS_reg_48_0_inst : DFFR_X1 port map( D => n7884, CK => CLK, RN => 
                           n3082, Q => n10117, QN => n1647);
   REGISTERS_reg_55_31_inst : DFFR_X1 port map( D => n8077, CK => CLK, RN => 
                           n3056, Q => n10118, QN => n1840);
   REGISTERS_reg_55_30_inst : DFFR_X1 port map( D => n8078, CK => CLK, RN => 
                           n3056, Q => n10119, QN => n1841);
   REGISTERS_reg_55_29_inst : DFFR_X1 port map( D => n8079, CK => CLK, RN => 
                           n3056, Q => n10120, QN => n1842);
   REGISTERS_reg_55_28_inst : DFFR_X1 port map( D => n8080, CK => CLK, RN => 
                           n3056, Q => n10121, QN => n1843);
   REGISTERS_reg_55_27_inst : DFFR_X1 port map( D => n8081, CK => CLK, RN => 
                           n3056, Q => n10122, QN => n1844);
   REGISTERS_reg_55_26_inst : DFFR_X1 port map( D => n8082, CK => CLK, RN => 
                           n3056, Q => n10123, QN => n1845);
   REGISTERS_reg_55_25_inst : DFFR_X1 port map( D => n8083, CK => CLK, RN => 
                           n3056, Q => n10124, QN => n1846);
   REGISTERS_reg_55_24_inst : DFFR_X1 port map( D => n8084, CK => CLK, RN => 
                           n3056, Q => n10125, QN => n1847);
   REGISTERS_reg_55_23_inst : DFFR_X1 port map( D => n8085, CK => CLK, RN => 
                           n3054, Q => n10126, QN => n1848);
   REGISTERS_reg_55_22_inst : DFFR_X1 port map( D => n8086, CK => CLK, RN => 
                           n3054, Q => n10127, QN => n1849);
   REGISTERS_reg_55_21_inst : DFFR_X1 port map( D => n8087, CK => CLK, RN => 
                           n3054, Q => n10128, QN => n1850);
   REGISTERS_reg_55_20_inst : DFFR_X1 port map( D => n8088, CK => CLK, RN => 
                           n3054, Q => n10129, QN => n1851);
   REGISTERS_reg_55_19_inst : DFFR_X1 port map( D => n8089, CK => CLK, RN => 
                           n3054, Q => n10130, QN => n1852);
   REGISTERS_reg_55_18_inst : DFFR_X1 port map( D => n8090, CK => CLK, RN => 
                           n3054, Q => n10131, QN => n1853);
   REGISTERS_reg_55_17_inst : DFFR_X1 port map( D => n8091, CK => CLK, RN => 
                           n3054, Q => n10132, QN => n1854);
   REGISTERS_reg_55_16_inst : DFFR_X1 port map( D => n8092, CK => CLK, RN => 
                           n3054, Q => n10133, QN => n1855);
   REGISTERS_reg_55_15_inst : DFFR_X1 port map( D => n8093, CK => CLK, RN => 
                           n3054, Q => n10134, QN => n1856);
   REGISTERS_reg_55_14_inst : DFFR_X1 port map( D => n8094, CK => CLK, RN => 
                           n3054, Q => n10135, QN => n1857);
   REGISTERS_reg_55_13_inst : DFFR_X1 port map( D => n8095, CK => CLK, RN => 
                           n3054, Q => n10136, QN => n1858);
   REGISTERS_reg_55_12_inst : DFFR_X1 port map( D => n8096, CK => CLK, RN => 
                           n3054, Q => n10137, QN => n1859);
   REGISTERS_reg_55_11_inst : DFFR_X1 port map( D => n8097, CK => CLK, RN => 
                           n3052, Q => n10138, QN => n1860);
   REGISTERS_reg_55_10_inst : DFFR_X1 port map( D => n8098, CK => CLK, RN => 
                           n3052, Q => n10139, QN => n1861);
   REGISTERS_reg_55_9_inst : DFFR_X1 port map( D => n8099, CK => CLK, RN => 
                           n3052, Q => n10140, QN => n1862);
   REGISTERS_reg_55_8_inst : DFFR_X1 port map( D => n8100, CK => CLK, RN => 
                           n3052, Q => n10141, QN => n1863);
   REGISTERS_reg_55_7_inst : DFFR_X1 port map( D => n8101, CK => CLK, RN => 
                           n3052, Q => n10142, QN => n1864);
   REGISTERS_reg_55_6_inst : DFFR_X1 port map( D => n8102, CK => CLK, RN => 
                           n3052, Q => n10143, QN => n1865);
   REGISTERS_reg_55_5_inst : DFFR_X1 port map( D => n8103, CK => CLK, RN => 
                           n3052, Q => n10144, QN => n1866);
   REGISTERS_reg_55_4_inst : DFFR_X1 port map( D => n8104, CK => CLK, RN => 
                           n3052, Q => n10145, QN => n1867);
   REGISTERS_reg_55_3_inst : DFFR_X1 port map( D => n8105, CK => CLK, RN => 
                           n3052, Q => n10146, QN => n1868);
   REGISTERS_reg_55_2_inst : DFFR_X1 port map( D => n8106, CK => CLK, RN => 
                           n3052, Q => n10147, QN => n1869);
   REGISTERS_reg_55_1_inst : DFFR_X1 port map( D => n8107, CK => CLK, RN => 
                           n3052, Q => n10148, QN => n1870);
   REGISTERS_reg_55_0_inst : DFFR_X1 port map( D => n8108, CK => CLK, RN => 
                           n3052, Q => n10149, QN => n1871);
   REGISTERS_reg_56_31_inst : DFFR_X1 port map( D => n8109, CK => CLK, RN => 
                           n3051, Q => n10150, QN => n1872);
   REGISTERS_reg_56_30_inst : DFFR_X1 port map( D => n8110, CK => CLK, RN => 
                           n3051, Q => n10151, QN => n1873);
   REGISTERS_reg_56_29_inst : DFFR_X1 port map( D => n8111, CK => CLK, RN => 
                           n3051, Q => n10152, QN => n1874);
   REGISTERS_reg_56_28_inst : DFFR_X1 port map( D => n8112, CK => CLK, RN => 
                           n3051, Q => n10153, QN => n1875);
   REGISTERS_reg_56_27_inst : DFFR_X1 port map( D => n8113, CK => CLK, RN => 
                           n3051, Q => n10154, QN => n1876);
   REGISTERS_reg_56_26_inst : DFFR_X1 port map( D => n8114, CK => CLK, RN => 
                           n3051, Q => n10155, QN => n1877);
   REGISTERS_reg_56_25_inst : DFFR_X1 port map( D => n8115, CK => CLK, RN => 
                           n3051, Q => n10156, QN => n1878);
   REGISTERS_reg_56_24_inst : DFFR_X1 port map( D => n8116, CK => CLK, RN => 
                           n3051, Q => n10157, QN => n1879);
   REGISTERS_reg_56_23_inst : DFFR_X1 port map( D => n8117, CK => CLK, RN => 
                           n3051, Q => n10158, QN => n1880);
   REGISTERS_reg_56_22_inst : DFFR_X1 port map( D => n8118, CK => CLK, RN => 
                           n3051, Q => n10159, QN => n1881);
   REGISTERS_reg_56_21_inst : DFFR_X1 port map( D => n8119, CK => CLK, RN => 
                           n3051, Q => n10160, QN => n1882);
   REGISTERS_reg_56_20_inst : DFFR_X1 port map( D => n8120, CK => CLK, RN => 
                           n3051, Q => n10161, QN => n1883);
   REGISTERS_reg_56_19_inst : DFFR_X1 port map( D => n8121, CK => CLK, RN => 
                           n3049, Q => n10162, QN => n1884);
   REGISTERS_reg_56_18_inst : DFFR_X1 port map( D => n8122, CK => CLK, RN => 
                           n3049, Q => n10163, QN => n1885);
   REGISTERS_reg_56_17_inst : DFFR_X1 port map( D => n8123, CK => CLK, RN => 
                           n3049, Q => n10164, QN => n1886);
   REGISTERS_reg_56_16_inst : DFFR_X1 port map( D => n8124, CK => CLK, RN => 
                           n3049, Q => n10165, QN => n1887);
   REGISTERS_reg_56_15_inst : DFFR_X1 port map( D => n8125, CK => CLK, RN => 
                           n3049, Q => n10166, QN => n1888);
   REGISTERS_reg_56_14_inst : DFFR_X1 port map( D => n8126, CK => CLK, RN => 
                           n3049, Q => n10167, QN => n1889);
   REGISTERS_reg_56_13_inst : DFFR_X1 port map( D => n8127, CK => CLK, RN => 
                           n3049, Q => n10168, QN => n1890);
   REGISTERS_reg_56_12_inst : DFFR_X1 port map( D => n8128, CK => CLK, RN => 
                           n3049, Q => n10169, QN => n1891);
   REGISTERS_reg_56_11_inst : DFFR_X1 port map( D => n8129, CK => CLK, RN => 
                           n3049, Q => n10170, QN => n1892);
   REGISTERS_reg_56_10_inst : DFFR_X1 port map( D => n8130, CK => CLK, RN => 
                           n3049, Q => n10171, QN => n1893);
   REGISTERS_reg_56_9_inst : DFFR_X1 port map( D => n8131, CK => CLK, RN => 
                           n3049, Q => n10172, QN => n1894);
   REGISTERS_reg_56_8_inst : DFFR_X1 port map( D => n8132, CK => CLK, RN => 
                           n3049, Q => n10173, QN => n1895);
   REGISTERS_reg_56_7_inst : DFFR_X1 port map( D => n8133, CK => CLK, RN => 
                           n3047, Q => n10174, QN => n1896);
   REGISTERS_reg_56_6_inst : DFFR_X1 port map( D => n8134, CK => CLK, RN => 
                           n3047, Q => n10175, QN => n1897);
   REGISTERS_reg_56_5_inst : DFFR_X1 port map( D => n8135, CK => CLK, RN => 
                           n3047, Q => n10176, QN => n1898);
   REGISTERS_reg_56_4_inst : DFFR_X1 port map( D => n8136, CK => CLK, RN => 
                           n3047, Q => n10177, QN => n1899);
   REGISTERS_reg_56_3_inst : DFFR_X1 port map( D => n8137, CK => CLK, RN => 
                           n3047, Q => n10178, QN => n1900);
   REGISTERS_reg_56_2_inst : DFFR_X1 port map( D => n8138, CK => CLK, RN => 
                           n3047, Q => n10179, QN => n1901);
   REGISTERS_reg_56_1_inst : DFFR_X1 port map( D => n8139, CK => CLK, RN => 
                           n3047, Q => n10180, QN => n1902);
   REGISTERS_reg_56_0_inst : DFFR_X1 port map( D => n8140, CK => CLK, RN => 
                           n3047, Q => n10181, QN => n1903);
   REGISTERS_reg_57_31_inst : DFFR_X1 port map( D => n8141, CK => CLK, RN => 
                           n3047, Q => n10182, QN => n1904);
   REGISTERS_reg_57_30_inst : DFFR_X1 port map( D => n8142, CK => CLK, RN => 
                           n3047, Q => n10183, QN => n1905);
   REGISTERS_reg_57_29_inst : DFFR_X1 port map( D => n8143, CK => CLK, RN => 
                           n3047, Q => n10184, QN => n1906);
   REGISTERS_reg_57_28_inst : DFFR_X1 port map( D => n8144, CK => CLK, RN => 
                           n3047, Q => n10185, QN => n1907);
   REGISTERS_reg_57_27_inst : DFFR_X1 port map( D => n8145, CK => CLK, RN => 
                           n3046, Q => n10186, QN => n1908);
   REGISTERS_reg_57_26_inst : DFFR_X1 port map( D => n8146, CK => CLK, RN => 
                           n3046, Q => n10187, QN => n1909);
   REGISTERS_reg_57_25_inst : DFFR_X1 port map( D => n8147, CK => CLK, RN => 
                           n3046, Q => n10188, QN => n1910);
   REGISTERS_reg_57_24_inst : DFFR_X1 port map( D => n8148, CK => CLK, RN => 
                           n3046, Q => n10189, QN => n1911);
   REGISTERS_reg_57_23_inst : DFFR_X1 port map( D => n8149, CK => CLK, RN => 
                           n3046, Q => n10190, QN => n1912);
   REGISTERS_reg_57_22_inst : DFFR_X1 port map( D => n8150, CK => CLK, RN => 
                           n3046, Q => n10191, QN => n1913);
   REGISTERS_reg_57_21_inst : DFFR_X1 port map( D => n8151, CK => CLK, RN => 
                           n3046, Q => n10192, QN => n1914);
   REGISTERS_reg_57_20_inst : DFFR_X1 port map( D => n8152, CK => CLK, RN => 
                           n3046, Q => n10193, QN => n1915);
   REGISTERS_reg_57_19_inst : DFFR_X1 port map( D => n8153, CK => CLK, RN => 
                           n3046, Q => n10194, QN => n1916);
   REGISTERS_reg_57_18_inst : DFFR_X1 port map( D => n8154, CK => CLK, RN => 
                           n3046, Q => n10195, QN => n1917);
   REGISTERS_reg_57_17_inst : DFFR_X1 port map( D => n8155, CK => CLK, RN => 
                           n3046, Q => n10196, QN => n1918);
   REGISTERS_reg_57_16_inst : DFFR_X1 port map( D => n8156, CK => CLK, RN => 
                           n3046, Q => n10197, QN => n1919);
   REGISTERS_reg_57_15_inst : DFFR_X1 port map( D => n8157, CK => CLK, RN => 
                           n3044, Q => n10198, QN => n1920);
   REGISTERS_reg_57_14_inst : DFFR_X1 port map( D => n8158, CK => CLK, RN => 
                           n3044, Q => n10199, QN => n1921);
   REGISTERS_reg_57_13_inst : DFFR_X1 port map( D => n8159, CK => CLK, RN => 
                           n3044, Q => n10200, QN => n1922);
   REGISTERS_reg_57_12_inst : DFFR_X1 port map( D => n8160, CK => CLK, RN => 
                           n3044, Q => n10201, QN => n1923);
   REGISTERS_reg_57_11_inst : DFFR_X1 port map( D => n8161, CK => CLK, RN => 
                           n3044, Q => n10202, QN => n1924);
   REGISTERS_reg_57_10_inst : DFFR_X1 port map( D => n8162, CK => CLK, RN => 
                           n3044, Q => n10203, QN => n1925);
   REGISTERS_reg_57_9_inst : DFFR_X1 port map( D => n8163, CK => CLK, RN => 
                           n3044, Q => n10204, QN => n1926);
   REGISTERS_reg_57_8_inst : DFFR_X1 port map( D => n8164, CK => CLK, RN => 
                           n3044, Q => n10205, QN => n1927);
   REGISTERS_reg_57_7_inst : DFFR_X1 port map( D => n8165, CK => CLK, RN => 
                           n3044, Q => n10206, QN => n1928);
   REGISTERS_reg_57_6_inst : DFFR_X1 port map( D => n8166, CK => CLK, RN => 
                           n3044, Q => n10207, QN => n1929);
   REGISTERS_reg_57_5_inst : DFFR_X1 port map( D => n8167, CK => CLK, RN => 
                           n3044, Q => n10208, QN => n1930);
   REGISTERS_reg_57_4_inst : DFFR_X1 port map( D => n8168, CK => CLK, RN => 
                           n3044, Q => n10209, QN => n1931);
   REGISTERS_reg_57_3_inst : DFFR_X1 port map( D => n8169, CK => CLK, RN => 
                           n3042, Q => n10210, QN => n1932);
   REGISTERS_reg_57_2_inst : DFFR_X1 port map( D => n8170, CK => CLK, RN => 
                           n3042, Q => n10211, QN => n1933);
   REGISTERS_reg_57_1_inst : DFFR_X1 port map( D => n8171, CK => CLK, RN => 
                           n3042, Q => n10212, QN => n1934);
   REGISTERS_reg_57_0_inst : DFFR_X1 port map( D => n8172, CK => CLK, RN => 
                           n3042, Q => n10213, QN => n1935);
   REGISTERS_reg_58_31_inst : DFFR_X1 port map( D => n8173, CK => CLK, RN => 
                           n3042, Q => n10214, QN => n1936);
   REGISTERS_reg_58_30_inst : DFFR_X1 port map( D => n8174, CK => CLK, RN => 
                           n3042, Q => n10215, QN => n1937);
   REGISTERS_reg_58_29_inst : DFFR_X1 port map( D => n8175, CK => CLK, RN => 
                           n3042, Q => n10216, QN => n1938);
   REGISTERS_reg_58_28_inst : DFFR_X1 port map( D => n8176, CK => CLK, RN => 
                           n3042, Q => n10217, QN => n1939);
   REGISTERS_reg_58_27_inst : DFFR_X1 port map( D => n8177, CK => CLK, RN => 
                           n3042, Q => n10218, QN => n1940);
   REGISTERS_reg_58_26_inst : DFFR_X1 port map( D => n8178, CK => CLK, RN => 
                           n3042, Q => n10219, QN => n1941);
   REGISTERS_reg_58_25_inst : DFFR_X1 port map( D => n8179, CK => CLK, RN => 
                           n3042, Q => n10220, QN => n1942);
   REGISTERS_reg_58_24_inst : DFFR_X1 port map( D => n8180, CK => CLK, RN => 
                           n3042, Q => n10221, QN => n1943);
   REGISTERS_reg_58_23_inst : DFFR_X1 port map( D => n8181, CK => CLK, RN => 
                           n3041, Q => n10222, QN => n1944);
   REGISTERS_reg_58_22_inst : DFFR_X1 port map( D => n8182, CK => CLK, RN => 
                           n3041, Q => n10223, QN => n1945);
   REGISTERS_reg_58_21_inst : DFFR_X1 port map( D => n8183, CK => CLK, RN => 
                           n3041, Q => n10224, QN => n1946);
   REGISTERS_reg_58_20_inst : DFFR_X1 port map( D => n8184, CK => CLK, RN => 
                           n3041, Q => n10225, QN => n1947);
   REGISTERS_reg_58_19_inst : DFFR_X1 port map( D => n8185, CK => CLK, RN => 
                           n3041, Q => n10226, QN => n1948);
   REGISTERS_reg_58_18_inst : DFFR_X1 port map( D => n8186, CK => CLK, RN => 
                           n3041, Q => n10227, QN => n1949);
   REGISTERS_reg_58_17_inst : DFFR_X1 port map( D => n8187, CK => CLK, RN => 
                           n3041, Q => n10228, QN => n1950);
   REGISTERS_reg_58_16_inst : DFFR_X1 port map( D => n8188, CK => CLK, RN => 
                           n3041, Q => n10229, QN => n1951);
   REGISTERS_reg_58_15_inst : DFFR_X1 port map( D => n8189, CK => CLK, RN => 
                           n3041, Q => n10230, QN => n1952);
   REGISTERS_reg_58_14_inst : DFFR_X1 port map( D => n8190, CK => CLK, RN => 
                           n3041, Q => n10231, QN => n1953);
   REGISTERS_reg_58_13_inst : DFFR_X1 port map( D => n8191, CK => CLK, RN => 
                           n3041, Q => n10232, QN => n1954);
   REGISTERS_reg_58_12_inst : DFFR_X1 port map( D => n8192, CK => CLK, RN => 
                           n3041, Q => n10233, QN => n1955);
   REGISTERS_reg_58_11_inst : DFFR_X1 port map( D => n8193, CK => CLK, RN => 
                           n3039, Q => n10234, QN => n1956);
   REGISTERS_reg_58_10_inst : DFFR_X1 port map( D => n8194, CK => CLK, RN => 
                           n3039, Q => n10235, QN => n1957);
   REGISTERS_reg_58_9_inst : DFFR_X1 port map( D => n8195, CK => CLK, RN => 
                           n3039, Q => n10236, QN => n1958);
   REGISTERS_reg_58_8_inst : DFFR_X1 port map( D => n8196, CK => CLK, RN => 
                           n3039, Q => n10237, QN => n1959);
   REGISTERS_reg_58_7_inst : DFFR_X1 port map( D => n8197, CK => CLK, RN => 
                           n3039, Q => n10238, QN => n1960);
   REGISTERS_reg_58_6_inst : DFFR_X1 port map( D => n8198, CK => CLK, RN => 
                           n3039, Q => n10239, QN => n1961);
   REGISTERS_reg_58_5_inst : DFFR_X1 port map( D => n8199, CK => CLK, RN => 
                           n3039, Q => n10240, QN => n1962);
   REGISTERS_reg_58_4_inst : DFFR_X1 port map( D => n8200, CK => CLK, RN => 
                           n3039, Q => n10241, QN => n1963);
   REGISTERS_reg_58_3_inst : DFFR_X1 port map( D => n8201, CK => CLK, RN => 
                           n3039, Q => n10242, QN => n1964);
   REGISTERS_reg_58_2_inst : DFFR_X1 port map( D => n8202, CK => CLK, RN => 
                           n3039, Q => n10243, QN => n1965);
   REGISTERS_reg_58_1_inst : DFFR_X1 port map( D => n8203, CK => CLK, RN => 
                           n3039, Q => n10244, QN => n1966);
   REGISTERS_reg_58_0_inst : DFFR_X1 port map( D => n8204, CK => CLK, RN => 
                           n3039, Q => n10245, QN => n1967);
   REGISTERS_reg_59_31_inst : DFFR_X1 port map( D => n8205, CK => CLK, RN => 
                           n3037, Q => n10246, QN => n1968);
   REGISTERS_reg_59_30_inst : DFFR_X1 port map( D => n8206, CK => CLK, RN => 
                           n3037, Q => n10247, QN => n1969);
   REGISTERS_reg_59_29_inst : DFFR_X1 port map( D => n8207, CK => CLK, RN => 
                           n3037, Q => n10248, QN => n1970);
   REGISTERS_reg_59_28_inst : DFFR_X1 port map( D => n8208, CK => CLK, RN => 
                           n3037, Q => n10249, QN => n1971);
   REGISTERS_reg_59_27_inst : DFFR_X1 port map( D => n8209, CK => CLK, RN => 
                           n3037, Q => n10250, QN => n1972);
   REGISTERS_reg_59_26_inst : DFFR_X1 port map( D => n8210, CK => CLK, RN => 
                           n3037, Q => n10251, QN => n1973);
   REGISTERS_reg_59_25_inst : DFFR_X1 port map( D => n8211, CK => CLK, RN => 
                           n3037, Q => n10252, QN => n1974);
   REGISTERS_reg_59_24_inst : DFFR_X1 port map( D => n8212, CK => CLK, RN => 
                           n3037, Q => n10253, QN => n1975);
   REGISTERS_reg_59_23_inst : DFFR_X1 port map( D => n8213, CK => CLK, RN => 
                           n3037, Q => n10254, QN => n1976);
   REGISTERS_reg_59_22_inst : DFFR_X1 port map( D => n8214, CK => CLK, RN => 
                           n3037, Q => n10255, QN => n1977);
   REGISTERS_reg_59_21_inst : DFFR_X1 port map( D => n8215, CK => CLK, RN => 
                           n3037, Q => n10256, QN => n1978);
   REGISTERS_reg_59_20_inst : DFFR_X1 port map( D => n8216, CK => CLK, RN => 
                           n3037, Q => n10257, QN => n1979);
   REGISTERS_reg_59_19_inst : DFFR_X1 port map( D => n8217, CK => CLK, RN => 
                           n3036, Q => n10258, QN => n1980);
   REGISTERS_reg_59_18_inst : DFFR_X1 port map( D => n8218, CK => CLK, RN => 
                           n3036, Q => n10259, QN => n1981);
   REGISTERS_reg_59_17_inst : DFFR_X1 port map( D => n8219, CK => CLK, RN => 
                           n3036, Q => n10260, QN => n1982);
   REGISTERS_reg_59_16_inst : DFFR_X1 port map( D => n8220, CK => CLK, RN => 
                           n3036, Q => n10261, QN => n1983);
   REGISTERS_reg_59_15_inst : DFFR_X1 port map( D => n8221, CK => CLK, RN => 
                           n3036, Q => n10262, QN => n1984);
   REGISTERS_reg_59_14_inst : DFFR_X1 port map( D => n8222, CK => CLK, RN => 
                           n3036, Q => n10263, QN => n1985);
   REGISTERS_reg_59_13_inst : DFFR_X1 port map( D => n8223, CK => CLK, RN => 
                           n3036, Q => n10264, QN => n1986);
   REGISTERS_reg_59_12_inst : DFFR_X1 port map( D => n8224, CK => CLK, RN => 
                           n3036, Q => n10265, QN => n1987);
   REGISTERS_reg_59_11_inst : DFFR_X1 port map( D => n8225, CK => CLK, RN => 
                           n3036, Q => n10266, QN => n1988);
   REGISTERS_reg_59_10_inst : DFFR_X1 port map( D => n8226, CK => CLK, RN => 
                           n3036, Q => n10267, QN => n1989);
   REGISTERS_reg_59_9_inst : DFFR_X1 port map( D => n8227, CK => CLK, RN => 
                           n3036, Q => n10268, QN => n1990);
   REGISTERS_reg_59_8_inst : DFFR_X1 port map( D => n8228, CK => CLK, RN => 
                           n3036, Q => n10269, QN => n1991);
   REGISTERS_reg_59_7_inst : DFFR_X1 port map( D => n8229, CK => CLK, RN => 
                           n3034, Q => n10270, QN => n1992);
   REGISTERS_reg_59_6_inst : DFFR_X1 port map( D => n8230, CK => CLK, RN => 
                           n3034, Q => n10271, QN => n1993);
   REGISTERS_reg_59_5_inst : DFFR_X1 port map( D => n8231, CK => CLK, RN => 
                           n3034, Q => n10272, QN => n1994);
   REGISTERS_reg_59_4_inst : DFFR_X1 port map( D => n8232, CK => CLK, RN => 
                           n3034, Q => n10273, QN => n1995);
   REGISTERS_reg_59_3_inst : DFFR_X1 port map( D => n8233, CK => CLK, RN => 
                           n3034, Q => n10274, QN => n1996);
   REGISTERS_reg_59_2_inst : DFFR_X1 port map( D => n8234, CK => CLK, RN => 
                           n3034, Q => n10275, QN => n1997);
   REGISTERS_reg_59_1_inst : DFFR_X1 port map( D => n8235, CK => CLK, RN => 
                           n3034, Q => n10276, QN => n1998);
   REGISTERS_reg_59_0_inst : DFFR_X1 port map( D => n8236, CK => CLK, RN => 
                           n3034, Q => n10277, QN => n1999);
   REGISTERS_reg_60_31_inst : DFFR_X1 port map( D => n8237, CK => CLK, RN => 
                           n3034, Q => n10278, QN => n2000);
   REGISTERS_reg_60_30_inst : DFFR_X1 port map( D => n8238, CK => CLK, RN => 
                           n3034, Q => n10279, QN => n2001);
   REGISTERS_reg_60_29_inst : DFFR_X1 port map( D => n8239, CK => CLK, RN => 
                           n3034, Q => n10280, QN => n2002);
   REGISTERS_reg_60_28_inst : DFFR_X1 port map( D => n8240, CK => CLK, RN => 
                           n3034, Q => n10281, QN => n2003);
   REGISTERS_reg_60_27_inst : DFFR_X1 port map( D => n8241, CK => CLK, RN => 
                           n3032, Q => n10282, QN => n2004);
   REGISTERS_reg_60_26_inst : DFFR_X1 port map( D => n8242, CK => CLK, RN => 
                           n3032, Q => n10283, QN => n2005);
   REGISTERS_reg_60_25_inst : DFFR_X1 port map( D => n8243, CK => CLK, RN => 
                           n3032, Q => n10284, QN => n2006);
   REGISTERS_reg_60_24_inst : DFFR_X1 port map( D => n8244, CK => CLK, RN => 
                           n3032, Q => n10285, QN => n2007);
   REGISTERS_reg_60_23_inst : DFFR_X1 port map( D => n8245, CK => CLK, RN => 
                           n3032, Q => n10286, QN => n2008);
   REGISTERS_reg_60_22_inst : DFFR_X1 port map( D => n8246, CK => CLK, RN => 
                           n3032, Q => n10287, QN => n2009);
   REGISTERS_reg_60_21_inst : DFFR_X1 port map( D => n8247, CK => CLK, RN => 
                           n3032, Q => n10288, QN => n2010);
   REGISTERS_reg_60_20_inst : DFFR_X1 port map( D => n8248, CK => CLK, RN => 
                           n3032, Q => n10289, QN => n2011);
   REGISTERS_reg_60_19_inst : DFFR_X1 port map( D => n8249, CK => CLK, RN => 
                           n3032, Q => n10290, QN => n2012);
   REGISTERS_reg_60_18_inst : DFFR_X1 port map( D => n8250, CK => CLK, RN => 
                           n3032, Q => n10291, QN => n2013);
   REGISTERS_reg_60_17_inst : DFFR_X1 port map( D => n8251, CK => CLK, RN => 
                           n3032, Q => n10292, QN => n2014);
   REGISTERS_reg_60_16_inst : DFFR_X1 port map( D => n8252, CK => CLK, RN => 
                           n3032, Q => n10293, QN => n2015);
   REGISTERS_reg_60_15_inst : DFFR_X1 port map( D => n8253, CK => CLK, RN => 
                           n3031, Q => n10294, QN => n2016);
   REGISTERS_reg_60_14_inst : DFFR_X1 port map( D => n8254, CK => CLK, RN => 
                           n3031, Q => n10295, QN => n2017);
   REGISTERS_reg_60_13_inst : DFFR_X1 port map( D => n8255, CK => CLK, RN => 
                           n3031, Q => n10296, QN => n2018);
   REGISTERS_reg_60_12_inst : DFFR_X1 port map( D => n8256, CK => CLK, RN => 
                           n3031, Q => n10297, QN => n2019);
   REGISTERS_reg_60_11_inst : DFFR_X1 port map( D => n8257, CK => CLK, RN => 
                           n3031, Q => n10298, QN => n2020);
   REGISTERS_reg_60_10_inst : DFFR_X1 port map( D => n8258, CK => CLK, RN => 
                           n3031, Q => n10299, QN => n2021);
   REGISTERS_reg_60_9_inst : DFFR_X1 port map( D => n8259, CK => CLK, RN => 
                           n3031, Q => n10300, QN => n2022);
   REGISTERS_reg_60_8_inst : DFFR_X1 port map( D => n8260, CK => CLK, RN => 
                           n3031, Q => n10301, QN => n2023);
   REGISTERS_reg_60_7_inst : DFFR_X1 port map( D => n8261, CK => CLK, RN => 
                           n3031, Q => n10302, QN => n2024);
   REGISTERS_reg_60_6_inst : DFFR_X1 port map( D => n8262, CK => CLK, RN => 
                           n3031, Q => n10303, QN => n2025);
   REGISTERS_reg_60_5_inst : DFFR_X1 port map( D => n8263, CK => CLK, RN => 
                           n3031, Q => n10304, QN => n2026);
   REGISTERS_reg_60_4_inst : DFFR_X1 port map( D => n8264, CK => CLK, RN => 
                           n3031, Q => n10305, QN => n2027);
   REGISTERS_reg_60_3_inst : DFFR_X1 port map( D => n8265, CK => CLK, RN => 
                           n3028, Q => n10306, QN => n2028);
   REGISTERS_reg_60_2_inst : DFFR_X1 port map( D => n8266, CK => CLK, RN => 
                           n3028, Q => n10307, QN => n2029);
   REGISTERS_reg_60_1_inst : DFFR_X1 port map( D => n8267, CK => CLK, RN => 
                           n3028, Q => n10308, QN => n2030);
   REGISTERS_reg_60_0_inst : DFFR_X1 port map( D => n8268, CK => CLK, RN => 
                           n3028, Q => n10309, QN => n2031);
   REGISTERS_reg_61_31_inst : DFFR_X1 port map( D => n8269, CK => CLK, RN => 
                           n3028, Q => n10310, QN => n2032);
   REGISTERS_reg_61_30_inst : DFFR_X1 port map( D => n8270, CK => CLK, RN => 
                           n3028, Q => n10311, QN => n2033);
   REGISTERS_reg_61_29_inst : DFFR_X1 port map( D => n8271, CK => CLK, RN => 
                           n3028, Q => n10312, QN => n2034);
   REGISTERS_reg_61_28_inst : DFFR_X1 port map( D => n8272, CK => CLK, RN => 
                           n3028, Q => n10313, QN => n2035);
   REGISTERS_reg_61_27_inst : DFFR_X1 port map( D => n8273, CK => CLK, RN => 
                           n3028, Q => n10314, QN => n2036);
   REGISTERS_reg_61_26_inst : DFFR_X1 port map( D => n8274, CK => CLK, RN => 
                           n3028, Q => n10315, QN => n2037);
   REGISTERS_reg_61_25_inst : DFFR_X1 port map( D => n8275, CK => CLK, RN => 
                           n3028, Q => n10316, QN => n2038);
   REGISTERS_reg_61_24_inst : DFFR_X1 port map( D => n8276, CK => CLK, RN => 
                           n3028, Q => n10317, QN => n2039);
   REGISTERS_reg_61_23_inst : DFFR_X1 port map( D => n8277, CK => CLK, RN => 
                           n3027, Q => n10318, QN => n2040);
   REGISTERS_reg_61_22_inst : DFFR_X1 port map( D => n8278, CK => CLK, RN => 
                           n3027, Q => n10319, QN => n2041);
   REGISTERS_reg_61_21_inst : DFFR_X1 port map( D => n8279, CK => CLK, RN => 
                           n3027, Q => n10320, QN => n2042);
   REGISTERS_reg_61_20_inst : DFFR_X1 port map( D => n8280, CK => CLK, RN => 
                           n3027, Q => n10321, QN => n2043);
   REGISTERS_reg_61_19_inst : DFFR_X1 port map( D => n8281, CK => CLK, RN => 
                           n3027, Q => n10322, QN => n2044);
   REGISTERS_reg_61_18_inst : DFFR_X1 port map( D => n8282, CK => CLK, RN => 
                           n3027, Q => n10323, QN => n2045);
   REGISTERS_reg_61_17_inst : DFFR_X1 port map( D => n8283, CK => CLK, RN => 
                           n3027, Q => n10324, QN => n2046);
   REGISTERS_reg_61_16_inst : DFFR_X1 port map( D => n8284, CK => CLK, RN => 
                           n3027, Q => n10325, QN => n2047);
   REGISTERS_reg_61_15_inst : DFFR_X1 port map( D => n8285, CK => CLK, RN => 
                           n3027, Q => n10326, QN => n2048);
   REGISTERS_reg_61_14_inst : DFFR_X1 port map( D => n8286, CK => CLK, RN => 
                           n3027, Q => n10327, QN => n2049);
   REGISTERS_reg_61_13_inst : DFFR_X1 port map( D => n8287, CK => CLK, RN => 
                           n3027, Q => n10328, QN => n2050);
   REGISTERS_reg_61_12_inst : DFFR_X1 port map( D => n8288, CK => CLK, RN => 
                           n3027, Q => n10329, QN => n2051);
   REGISTERS_reg_61_11_inst : DFFR_X1 port map( D => n8289, CK => CLK, RN => 
                           n3026, Q => n10330, QN => n2052);
   REGISTERS_reg_61_10_inst : DFFR_X1 port map( D => n8290, CK => CLK, RN => 
                           n3026, Q => n10331, QN => n2053);
   REGISTERS_reg_61_9_inst : DFFR_X1 port map( D => n8291, CK => CLK, RN => 
                           n3026, Q => n10332, QN => n2054);
   REGISTERS_reg_61_8_inst : DFFR_X1 port map( D => n8292, CK => CLK, RN => 
                           n3026, Q => n10333, QN => n2055);
   REGISTERS_reg_61_7_inst : DFFR_X1 port map( D => n8293, CK => CLK, RN => 
                           n3026, Q => n10334, QN => n2056);
   REGISTERS_reg_61_6_inst : DFFR_X1 port map( D => n8294, CK => CLK, RN => 
                           n3026, Q => n10335, QN => n2057);
   REGISTERS_reg_61_5_inst : DFFR_X1 port map( D => n8295, CK => CLK, RN => 
                           n3026, Q => n10336, QN => n2058);
   REGISTERS_reg_61_4_inst : DFFR_X1 port map( D => n8296, CK => CLK, RN => 
                           n3026, Q => n10337, QN => n2059);
   REGISTERS_reg_61_3_inst : DFFR_X1 port map( D => n8297, CK => CLK, RN => 
                           n3026, Q => n10338, QN => n2060);
   REGISTERS_reg_61_2_inst : DFFR_X1 port map( D => n8298, CK => CLK, RN => 
                           n3026, Q => n10339, QN => n2061);
   REGISTERS_reg_61_1_inst : DFFR_X1 port map( D => n8299, CK => CLK, RN => 
                           n3026, Q => n10340, QN => n2062);
   REGISTERS_reg_61_0_inst : DFFR_X1 port map( D => n8300, CK => CLK, RN => 
                           n3026, Q => n10341, QN => n2063);
   REGISTERS_reg_62_31_inst : DFFR_X1 port map( D => n8301, CK => CLK, RN => 
                           n2994, Q => n10342, QN => n2064);
   REGISTERS_reg_62_30_inst : DFFR_X1 port map( D => n8302, CK => CLK, RN => 
                           n2992, Q => n10343, QN => n2065);
   REGISTERS_reg_62_29_inst : DFFR_X1 port map( D => n8303, CK => CLK, RN => 
                           n3004, Q => n10344, QN => n2066);
   REGISTERS_reg_62_28_inst : DFFR_X1 port map( D => n8304, CK => CLK, RN => 
                           n3005, Q => n10345, QN => n2067);
   REGISTERS_reg_62_27_inst : DFFR_X1 port map( D => n8305, CK => CLK, RN => 
                           n2993, Q => n10346, QN => n2068);
   REGISTERS_reg_62_26_inst : DFFR_X1 port map( D => n8306, CK => CLK, RN => 
                           n3001, Q => n10347, QN => n2069);
   REGISTERS_reg_62_25_inst : DFFR_X1 port map( D => n8307, CK => CLK, RN => 
                           n3002, Q => n10348, QN => n2070);
   REGISTERS_reg_62_24_inst : DFFR_X1 port map( D => n8308, CK => CLK, RN => 
                           n2999, Q => n10349, QN => n2071);
   REGISTERS_reg_62_23_inst : DFFR_X1 port map( D => n8309, CK => CLK, RN => 
                           n2995, Q => n10350, QN => n2072);
   REGISTERS_reg_62_22_inst : DFFR_X1 port map( D => n8310, CK => CLK, RN => 
                           n3003, Q => n10351, QN => n2073);
   REGISTERS_reg_62_21_inst : DFFR_X1 port map( D => n8311, CK => CLK, RN => 
                           n3000, Q => n10352, QN => n2074);
   REGISTERS_reg_62_20_inst : DFFR_X1 port map( D => n8312, CK => CLK, RN => 
                           n2991, Q => n10353, QN => n2075);
   REGISTERS_reg_62_19_inst : DFFR_X1 port map( D => n8313, CK => CLK, RN => 
                           n3025, Q => n10354, QN => n2076);
   REGISTERS_reg_62_18_inst : DFFR_X1 port map( D => n8314, CK => CLK, RN => 
                           n3025, Q => n10355, QN => n2077);
   REGISTERS_reg_62_17_inst : DFFR_X1 port map( D => n8315, CK => CLK, RN => 
                           n3025, Q => n10356, QN => n2078);
   REGISTERS_reg_62_16_inst : DFFR_X1 port map( D => n8316, CK => CLK, RN => 
                           n3025, Q => n10357, QN => n2079);
   REGISTERS_reg_62_15_inst : DFFR_X1 port map( D => n8317, CK => CLK, RN => 
                           n3025, Q => n10358, QN => n2080);
   REGISTERS_reg_62_14_inst : DFFR_X1 port map( D => n8318, CK => CLK, RN => 
                           n3025, Q => n10359, QN => n2081);
   REGISTERS_reg_62_13_inst : DFFR_X1 port map( D => n8319, CK => CLK, RN => 
                           n3025, Q => n10360, QN => n2082);
   REGISTERS_reg_62_12_inst : DFFR_X1 port map( D => n8320, CK => CLK, RN => 
                           n3025, Q => n10361, QN => n2083);
   REGISTERS_reg_62_11_inst : DFFR_X1 port map( D => n8321, CK => CLK, RN => 
                           n3025, Q => n10362, QN => n2084);
   REGISTERS_reg_62_10_inst : DFFR_X1 port map( D => n8322, CK => CLK, RN => 
                           n3025, Q => n10363, QN => n2085);
   REGISTERS_reg_62_9_inst : DFFR_X1 port map( D => n8323, CK => CLK, RN => 
                           n3025, Q => n10364, QN => n2086);
   REGISTERS_reg_62_8_inst : DFFR_X1 port map( D => n8324, CK => CLK, RN => 
                           n3025, Q => n10365, QN => n2087);
   REGISTERS_reg_62_7_inst : DFFR_X1 port map( D => n8325, CK => CLK, RN => 
                           n3024, Q => n10366, QN => n2088);
   REGISTERS_reg_62_6_inst : DFFR_X1 port map( D => n8326, CK => CLK, RN => 
                           n3024, Q => n10367, QN => n2089);
   REGISTERS_reg_62_5_inst : DFFR_X1 port map( D => n8327, CK => CLK, RN => 
                           n3024, Q => n10368, QN => n2090);
   REGISTERS_reg_62_4_inst : DFFR_X1 port map( D => n8328, CK => CLK, RN => 
                           n3024, Q => n10369, QN => n2091);
   REGISTERS_reg_62_3_inst : DFFR_X1 port map( D => n8329, CK => CLK, RN => 
                           n3024, Q => n10370, QN => n2092);
   REGISTERS_reg_62_2_inst : DFFR_X1 port map( D => n8330, CK => CLK, RN => 
                           n3024, Q => n10371, QN => n2093);
   REGISTERS_reg_62_1_inst : DFFR_X1 port map( D => n8331, CK => CLK, RN => 
                           n3024, Q => n10372, QN => n2094);
   REGISTERS_reg_62_0_inst : DFFR_X1 port map( D => n8332, CK => CLK, RN => 
                           n3024, Q => n10373, QN => n2095);
   REGISTERS_reg_63_31_inst : DFFR_X1 port map( D => n8333, CK => CLK, RN => 
                           n3024, Q => n10374, QN => n2096);
   REGISTERS_reg_63_30_inst : DFFR_X1 port map( D => n8334, CK => CLK, RN => 
                           n3024, Q => n10375, QN => n2097);
   REGISTERS_reg_63_29_inst : DFFR_X1 port map( D => n8335, CK => CLK, RN => 
                           n3024, Q => n10376, QN => n2098);
   REGISTERS_reg_63_28_inst : DFFR_X1 port map( D => n8336, CK => CLK, RN => 
                           n3024, Q => n10377, QN => n2099);
   REGISTERS_reg_63_27_inst : DFFR_X1 port map( D => n8337, CK => CLK, RN => 
                           n3023, Q => n10378, QN => n2100);
   REGISTERS_reg_63_26_inst : DFFR_X1 port map( D => n8338, CK => CLK, RN => 
                           n3023, Q => n10379, QN => n2101);
   REGISTERS_reg_63_25_inst : DFFR_X1 port map( D => n8339, CK => CLK, RN => 
                           n3023, Q => n10380, QN => n2102);
   REGISTERS_reg_63_24_inst : DFFR_X1 port map( D => n8340, CK => CLK, RN => 
                           n3023, Q => n10381, QN => n2103);
   REGISTERS_reg_63_23_inst : DFFR_X1 port map( D => n8341, CK => CLK, RN => 
                           n3023, Q => n10382, QN => n2104);
   REGISTERS_reg_63_22_inst : DFFR_X1 port map( D => n8342, CK => CLK, RN => 
                           n3023, Q => n10383, QN => n2105);
   REGISTERS_reg_63_21_inst : DFFR_X1 port map( D => n8343, CK => CLK, RN => 
                           n3023, Q => n10384, QN => n2106);
   REGISTERS_reg_63_20_inst : DFFR_X1 port map( D => n8344, CK => CLK, RN => 
                           n3023, Q => n10385, QN => n2107);
   REGISTERS_reg_63_19_inst : DFFR_X1 port map( D => n8345, CK => CLK, RN => 
                           n3023, Q => n10386, QN => n2108);
   REGISTERS_reg_63_18_inst : DFFR_X1 port map( D => n8346, CK => CLK, RN => 
                           n3023, Q => n10387, QN => n2109);
   REGISTERS_reg_63_17_inst : DFFR_X1 port map( D => n8347, CK => CLK, RN => 
                           n3023, Q => n10388, QN => n2110);
   REGISTERS_reg_63_16_inst : DFFR_X1 port map( D => n8348, CK => CLK, RN => 
                           n3023, Q => n10389, QN => n2111);
   REGISTERS_reg_63_15_inst : DFFR_X1 port map( D => n8349, CK => CLK, RN => 
                           n3022, Q => n10390, QN => n2112);
   REGISTERS_reg_63_14_inst : DFFR_X1 port map( D => n8350, CK => CLK, RN => 
                           n3022, Q => n10391, QN => n2113);
   REGISTERS_reg_63_13_inst : DFFR_X1 port map( D => n8351, CK => CLK, RN => 
                           n3022, Q => n10392, QN => n2114);
   REGISTERS_reg_63_12_inst : DFFR_X1 port map( D => n8352, CK => CLK, RN => 
                           n3022, Q => n10393, QN => n2115);
   REGISTERS_reg_63_11_inst : DFFR_X1 port map( D => n8353, CK => CLK, RN => 
                           n3022, Q => n10394, QN => n2116);
   REGISTERS_reg_63_10_inst : DFFR_X1 port map( D => n8354, CK => CLK, RN => 
                           n3022, Q => n10395, QN => n2117);
   REGISTERS_reg_63_9_inst : DFFR_X1 port map( D => n8355, CK => CLK, RN => 
                           n3022, Q => n10396, QN => n2118);
   REGISTERS_reg_63_8_inst : DFFR_X1 port map( D => n8356, CK => CLK, RN => 
                           n3022, Q => n10397, QN => n2119);
   REGISTERS_reg_63_7_inst : DFFR_X1 port map( D => n8357, CK => CLK, RN => 
                           n3022, Q => n10398, QN => n2120);
   REGISTERS_reg_63_6_inst : DFFR_X1 port map( D => n8358, CK => CLK, RN => 
                           n3022, Q => n10399, QN => n2121);
   REGISTERS_reg_63_5_inst : DFFR_X1 port map( D => n8359, CK => CLK, RN => 
                           n3022, Q => n10400, QN => n2122);
   REGISTERS_reg_63_4_inst : DFFR_X1 port map( D => n8360, CK => CLK, RN => 
                           n3022, Q => n10401, QN => n2123);
   REGISTERS_reg_63_3_inst : DFFR_X1 port map( D => n8361, CK => CLK, RN => 
                           n3021, Q => n10402, QN => n2124);
   REGISTERS_reg_63_2_inst : DFFR_X1 port map( D => n8362, CK => CLK, RN => 
                           n3021, Q => n10403, QN => n2125);
   REGISTERS_reg_63_1_inst : DFFR_X1 port map( D => n8363, CK => CLK, RN => 
                           n3021, Q => n10404, QN => n2126);
   REGISTERS_reg_63_0_inst : DFFR_X1 port map( D => n8364, CK => CLK, RN => 
                           n3021, Q => n10405, QN => n2127);
   REGISTERS_reg_64_31_inst : DFFR_X1 port map( D => n8365, CK => CLK, RN => 
                           n3021, Q => n10406, QN => n2128);
   REGISTERS_reg_64_30_inst : DFFR_X1 port map( D => n8366, CK => CLK, RN => 
                           n3021, Q => n10407, QN => n2129);
   REGISTERS_reg_64_29_inst : DFFR_X1 port map( D => n8367, CK => CLK, RN => 
                           n3021, Q => n10408, QN => n2130);
   REGISTERS_reg_64_28_inst : DFFR_X1 port map( D => n8368, CK => CLK, RN => 
                           n3021, Q => n10409, QN => n2131);
   REGISTERS_reg_64_27_inst : DFFR_X1 port map( D => n8369, CK => CLK, RN => 
                           n3021, Q => n10410, QN => n2132);
   REGISTERS_reg_64_26_inst : DFFR_X1 port map( D => n8370, CK => CLK, RN => 
                           n3021, Q => n10411, QN => n2133);
   REGISTERS_reg_64_25_inst : DFFR_X1 port map( D => n8371, CK => CLK, RN => 
                           n3021, Q => n10412, QN => n2134);
   REGISTERS_reg_64_24_inst : DFFR_X1 port map( D => n8372, CK => CLK, RN => 
                           n3021, Q => n10413, QN => n2135);
   REGISTERS_reg_64_23_inst : DFFR_X1 port map( D => n8373, CK => CLK, RN => 
                           n3020, Q => n10414, QN => n2136);
   REGISTERS_reg_64_22_inst : DFFR_X1 port map( D => n8374, CK => CLK, RN => 
                           n3020, Q => n10415, QN => n2137);
   REGISTERS_reg_64_21_inst : DFFR_X1 port map( D => n8375, CK => CLK, RN => 
                           n3020, Q => n10416, QN => n2138);
   REGISTERS_reg_64_20_inst : DFFR_X1 port map( D => n8376, CK => CLK, RN => 
                           n3020, Q => n10417, QN => n2139);
   REGISTERS_reg_64_19_inst : DFFR_X1 port map( D => n8377, CK => CLK, RN => 
                           n3020, Q => n10418, QN => n2140);
   REGISTERS_reg_64_18_inst : DFFR_X1 port map( D => n8378, CK => CLK, RN => 
                           n3020, Q => n10419, QN => n2141);
   REGISTERS_reg_64_17_inst : DFFR_X1 port map( D => n8379, CK => CLK, RN => 
                           n3020, Q => n10420, QN => n2142);
   REGISTERS_reg_64_16_inst : DFFR_X1 port map( D => n8380, CK => CLK, RN => 
                           n3020, Q => n10421, QN => n2143);
   REGISTERS_reg_64_15_inst : DFFR_X1 port map( D => n8381, CK => CLK, RN => 
                           n3020, Q => n10422, QN => n2144);
   REGISTERS_reg_64_14_inst : DFFR_X1 port map( D => n8382, CK => CLK, RN => 
                           n3020, Q => n10423, QN => n2145);
   REGISTERS_reg_64_13_inst : DFFR_X1 port map( D => n8383, CK => CLK, RN => 
                           n3020, Q => n10424, QN => n2146);
   REGISTERS_reg_64_12_inst : DFFR_X1 port map( D => n8384, CK => CLK, RN => 
                           n3020, Q => n10425, QN => n2147);
   REGISTERS_reg_64_11_inst : DFFR_X1 port map( D => n8385, CK => CLK, RN => 
                           n3019, Q => n10426, QN => n2148);
   REGISTERS_reg_64_10_inst : DFFR_X1 port map( D => n8386, CK => CLK, RN => 
                           n3019, Q => n10427, QN => n2149);
   REGISTERS_reg_64_9_inst : DFFR_X1 port map( D => n8387, CK => CLK, RN => 
                           n3019, Q => n10428, QN => n2150);
   REGISTERS_reg_64_8_inst : DFFR_X1 port map( D => n8388, CK => CLK, RN => 
                           n3019, Q => n10429, QN => n2151_port);
   REGISTERS_reg_64_7_inst : DFFR_X1 port map( D => n8389, CK => CLK, RN => 
                           n3019, Q => n10430, QN => n2152);
   REGISTERS_reg_64_6_inst : DFFR_X1 port map( D => n8390, CK => CLK, RN => 
                           n3019, Q => n10431, QN => n2153_port);
   REGISTERS_reg_64_5_inst : DFFR_X1 port map( D => n8391, CK => CLK, RN => 
                           n3019, Q => n10432, QN => n2154_port);
   REGISTERS_reg_64_4_inst : DFFR_X1 port map( D => n8392, CK => CLK, RN => 
                           n3019, Q => n10433, QN => n2155_port);
   REGISTERS_reg_64_3_inst : DFFR_X1 port map( D => n8393, CK => CLK, RN => 
                           n3019, Q => n10434, QN => n2156_port);
   REGISTERS_reg_64_2_inst : DFFR_X1 port map( D => n8394, CK => CLK, RN => 
                           n3019, Q => n10435, QN => n2157_port);
   REGISTERS_reg_64_1_inst : DFFR_X1 port map( D => n8395, CK => CLK, RN => 
                           n3019, Q => n10436, QN => n2158_port);
   REGISTERS_reg_64_0_inst : DFFR_X1 port map( D => n8396, CK => CLK, RN => 
                           n3019, Q => n10437, QN => n2159_port);
   REGISTERS_reg_65_31_inst : DFFR_X1 port map( D => n8397, CK => CLK, RN => 
                           n3018, Q => n10438, QN => n2160);
   REGISTERS_reg_65_30_inst : DFFR_X1 port map( D => n8398, CK => CLK, RN => 
                           n3018, Q => n10439, QN => n2161);
   REGISTERS_reg_65_29_inst : DFFR_X1 port map( D => n8399, CK => CLK, RN => 
                           n3018, Q => n10440, QN => n2162);
   REGISTERS_reg_65_28_inst : DFFR_X1 port map( D => n8400, CK => CLK, RN => 
                           n3018, Q => n10441, QN => n2163_port);
   REGISTERS_reg_65_27_inst : DFFR_X1 port map( D => n8401, CK => CLK, RN => 
                           n3018, Q => n10442, QN => n2164_port);
   REGISTERS_reg_65_26_inst : DFFR_X1 port map( D => n8402, CK => CLK, RN => 
                           n3018, Q => n10443, QN => n2165_port);
   REGISTERS_reg_65_25_inst : DFFR_X1 port map( D => n8403, CK => CLK, RN => 
                           n3018, Q => n10444, QN => n2166_port);
   REGISTERS_reg_65_24_inst : DFFR_X1 port map( D => n8404, CK => CLK, RN => 
                           n3018, Q => n10445, QN => n2167);
   REGISTERS_reg_65_23_inst : DFFR_X1 port map( D => n8405, CK => CLK, RN => 
                           n3018, Q => n10446, QN => n2168);
   REGISTERS_reg_65_22_inst : DFFR_X1 port map( D => n8406, CK => CLK, RN => 
                           n3018, Q => n10447, QN => n2169);
   REGISTERS_reg_65_21_inst : DFFR_X1 port map( D => n8407, CK => CLK, RN => 
                           n3018, Q => n10448, QN => n2170);
   REGISTERS_reg_65_20_inst : DFFR_X1 port map( D => n8408, CK => CLK, RN => 
                           n3018, Q => n10449, QN => n2171);
   REGISTERS_reg_65_19_inst : DFFR_X1 port map( D => n8409, CK => CLK, RN => 
                           n3017, Q => n10450, QN => n2172);
   REGISTERS_reg_65_18_inst : DFFR_X1 port map( D => n8410, CK => CLK, RN => 
                           n3017, Q => n10451, QN => n2173);
   REGISTERS_reg_65_17_inst : DFFR_X1 port map( D => n8411, CK => CLK, RN => 
                           n3017, Q => n10452, QN => n2174);
   REGISTERS_reg_65_16_inst : DFFR_X1 port map( D => n8412, CK => CLK, RN => 
                           n3017, Q => n10453, QN => n2175);
   REGISTERS_reg_65_15_inst : DFFR_X1 port map( D => n8413, CK => CLK, RN => 
                           n3017, Q => n10454, QN => n2176);
   REGISTERS_reg_65_14_inst : DFFR_X1 port map( D => n8414, CK => CLK, RN => 
                           n3017, Q => n10455, QN => n2177);
   REGISTERS_reg_65_13_inst : DFFR_X1 port map( D => n8415_port, CK => CLK, RN 
                           => n3017, Q => n10456, QN => n2178);
   REGISTERS_reg_65_12_inst : DFFR_X1 port map( D => n8416, CK => CLK, RN => 
                           n3017, Q => n10457, QN => n2179);
   REGISTERS_reg_65_11_inst : DFFR_X1 port map( D => n8417_port, CK => CLK, RN 
                           => n3017, Q => n10458, QN => n2180);
   REGISTERS_reg_65_10_inst : DFFR_X1 port map( D => n8418_port, CK => CLK, RN 
                           => n3017, Q => n10459, QN => n2181);
   REGISTERS_reg_65_9_inst : DFFR_X1 port map( D => n8419_port, CK => CLK, RN 
                           => n3017, Q => n10460, QN => n2182);
   REGISTERS_reg_65_8_inst : DFFR_X1 port map( D => n8420_port, CK => CLK, RN 
                           => n3017, Q => n10461, QN => n2183);
   REGISTERS_reg_65_7_inst : DFFR_X1 port map( D => n8421_port, CK => CLK, RN 
                           => n3016, Q => n10462, QN => n2184);
   REGISTERS_reg_65_6_inst : DFFR_X1 port map( D => n8422_port, CK => CLK, RN 
                           => n3016, Q => n10463, QN => n2185);
   REGISTERS_reg_65_5_inst : DFFR_X1 port map( D => n8423_port, CK => CLK, RN 
                           => n3016, Q => n10464, QN => n2186);
   REGISTERS_reg_65_4_inst : DFFR_X1 port map( D => n8424, CK => CLK, RN => 
                           n3016, Q => n10465, QN => n2187);
   REGISTERS_reg_65_3_inst : DFFR_X1 port map( D => n8425, CK => CLK, RN => 
                           n3016, Q => n10466, QN => n2188);
   REGISTERS_reg_65_2_inst : DFFR_X1 port map( D => n8426, CK => CLK, RN => 
                           n3016, Q => n10467, QN => n2189);
   REGISTERS_reg_65_1_inst : DFFR_X1 port map( D => n8427_port, CK => CLK, RN 
                           => n3016, Q => n10468, QN => n2190);
   REGISTERS_reg_65_0_inst : DFFR_X1 port map( D => n8428_port, CK => CLK, RN 
                           => n3016, Q => n10469, QN => n2191);
   REGISTERS_reg_66_31_inst : DFFR_X1 port map( D => n8429_port, CK => CLK, RN 
                           => n3016, Q => n10470, QN => n2192);
   REGISTERS_reg_66_30_inst : DFFR_X1 port map( D => n8430_port, CK => CLK, RN 
                           => n3016, Q => n10471, QN => n2193);
   REGISTERS_reg_66_29_inst : DFFR_X1 port map( D => n8431, CK => CLK, RN => 
                           n3016, Q => n10472, QN => n2194);
   REGISTERS_reg_66_28_inst : DFFR_X1 port map( D => n8432, CK => CLK, RN => 
                           n3016, Q => n10473, QN => n2195);
   REGISTERS_reg_66_27_inst : DFFR_X1 port map( D => n8433, CK => CLK, RN => 
                           n3015, Q => n10474, QN => n2196);
   REGISTERS_reg_66_26_inst : DFFR_X1 port map( D => n8434, CK => CLK, RN => 
                           n3015, Q => n10475, QN => n2197);
   REGISTERS_reg_66_25_inst : DFFR_X1 port map( D => n8435, CK => CLK, RN => 
                           n3015, Q => n10476, QN => n2198);
   REGISTERS_reg_66_24_inst : DFFR_X1 port map( D => n8436, CK => CLK, RN => 
                           n3015, Q => n10477, QN => n2199);
   REGISTERS_reg_66_23_inst : DFFR_X1 port map( D => n8437, CK => CLK, RN => 
                           n3015, Q => n10478, QN => n2200);
   REGISTERS_reg_66_22_inst : DFFR_X1 port map( D => n8438, CK => CLK, RN => 
                           n3015, Q => n10479, QN => n2201);
   REGISTERS_reg_66_21_inst : DFFR_X1 port map( D => n8439, CK => CLK, RN => 
                           n3015, Q => n10480, QN => n2202);
   REGISTERS_reg_66_20_inst : DFFR_X1 port map( D => n8440, CK => CLK, RN => 
                           n3015, Q => n10481, QN => n2203);
   REGISTERS_reg_66_19_inst : DFFR_X1 port map( D => n8441, CK => CLK, RN => 
                           n3015, Q => n10482, QN => n2204);
   REGISTERS_reg_66_18_inst : DFFR_X1 port map( D => n8442, CK => CLK, RN => 
                           n3015, Q => n10483, QN => n2205);
   REGISTERS_reg_66_17_inst : DFFR_X1 port map( D => n8443, CK => CLK, RN => 
                           n3015, Q => n10484, QN => n2206);
   REGISTERS_reg_66_16_inst : DFFR_X1 port map( D => n8444, CK => CLK, RN => 
                           n3015, Q => n10485, QN => n2207);
   REGISTERS_reg_66_15_inst : DFFR_X1 port map( D => n8445, CK => CLK, RN => 
                           n3014, Q => n10486, QN => n2208);
   REGISTERS_reg_66_14_inst : DFFR_X1 port map( D => n8446, CK => CLK, RN => 
                           n3014, Q => n10487, QN => n2209);
   REGISTERS_reg_66_13_inst : DFFR_X1 port map( D => n8447, CK => CLK, RN => 
                           n3014, Q => n10488, QN => n2210);
   REGISTERS_reg_66_12_inst : DFFR_X1 port map( D => n8448, CK => CLK, RN => 
                           n3014, Q => n10489, QN => n2211);
   REGISTERS_reg_66_11_inst : DFFR_X1 port map( D => n8449, CK => CLK, RN => 
                           n3014, Q => n10490, QN => n2212);
   REGISTERS_reg_66_10_inst : DFFR_X1 port map( D => n8450, CK => CLK, RN => 
                           n3014, Q => n10491, QN => n2213);
   REGISTERS_reg_66_9_inst : DFFR_X1 port map( D => n8451, CK => CLK, RN => 
                           n3014, Q => n10492, QN => n2214);
   REGISTERS_reg_66_8_inst : DFFR_X1 port map( D => n8452, CK => CLK, RN => 
                           n3014, Q => n10493, QN => n2215);
   REGISTERS_reg_66_7_inst : DFFR_X1 port map( D => n8453, CK => CLK, RN => 
                           n3014, Q => n10494, QN => n2216);
   REGISTERS_reg_66_6_inst : DFFR_X1 port map( D => n8454, CK => CLK, RN => 
                           n3014, Q => n10495, QN => n2217);
   REGISTERS_reg_66_5_inst : DFFR_X1 port map( D => n8455, CK => CLK, RN => 
                           n3014, Q => n10496, QN => n2218);
   REGISTERS_reg_66_4_inst : DFFR_X1 port map( D => n8456, CK => CLK, RN => 
                           n3014, Q => n10497, QN => n2219);
   REGISTERS_reg_66_3_inst : DFFR_X1 port map( D => n8457, CK => CLK, RN => 
                           n3013, Q => n10498, QN => n2220);
   REGISTERS_reg_66_2_inst : DFFR_X1 port map( D => n8458, CK => CLK, RN => 
                           n3013, Q => n10499, QN => n2221);
   REGISTERS_reg_66_1_inst : DFFR_X1 port map( D => n8459, CK => CLK, RN => 
                           n3013, Q => n10500, QN => n2222);
   REGISTERS_reg_66_0_inst : DFFR_X1 port map( D => n8460, CK => CLK, RN => 
                           n3013, Q => n10501, QN => n2223);
   REGISTERS_reg_67_31_inst : DFFR_X1 port map( D => n8461, CK => CLK, RN => 
                           n3013, Q => n10502, QN => n2224);
   REGISTERS_reg_67_30_inst : DFFR_X1 port map( D => n8462, CK => CLK, RN => 
                           n3013, Q => n10503, QN => n2225);
   REGISTERS_reg_67_29_inst : DFFR_X1 port map( D => n8463, CK => CLK, RN => 
                           n3013, Q => n10504, QN => n2226);
   REGISTERS_reg_67_28_inst : DFFR_X1 port map( D => n8464, CK => CLK, RN => 
                           n3013, Q => n10505, QN => n2227);
   REGISTERS_reg_67_27_inst : DFFR_X1 port map( D => n8465, CK => CLK, RN => 
                           n3013, Q => n10506, QN => n2228);
   REGISTERS_reg_67_26_inst : DFFR_X1 port map( D => n8466, CK => CLK, RN => 
                           n3013, Q => n10507, QN => n2229);
   REGISTERS_reg_67_25_inst : DFFR_X1 port map( D => n8467, CK => CLK, RN => 
                           n3013, Q => n10508, QN => n2230);
   REGISTERS_reg_67_24_inst : DFFR_X1 port map( D => n8468, CK => CLK, RN => 
                           n3013, Q => n10509, QN => n2231);
   REGISTERS_reg_67_23_inst : DFFR_X1 port map( D => n8469, CK => CLK, RN => 
                           n3012, Q => n10510, QN => n2232);
   REGISTERS_reg_67_22_inst : DFFR_X1 port map( D => n8470, CK => CLK, RN => 
                           n3012, Q => n10511, QN => n2233);
   REGISTERS_reg_67_21_inst : DFFR_X1 port map( D => n8471, CK => CLK, RN => 
                           n3012, Q => n10512, QN => n2234);
   REGISTERS_reg_67_20_inst : DFFR_X1 port map( D => n8472, CK => CLK, RN => 
                           n3012, Q => n10513, QN => n2235);
   REGISTERS_reg_67_19_inst : DFFR_X1 port map( D => n8473, CK => CLK, RN => 
                           n3012, Q => n10514, QN => n2236);
   REGISTERS_reg_67_18_inst : DFFR_X1 port map( D => n8474, CK => CLK, RN => 
                           n3012, Q => n10515, QN => n2237);
   REGISTERS_reg_67_17_inst : DFFR_X1 port map( D => n8475, CK => CLK, RN => 
                           n3012, Q => n10516, QN => n2238);
   REGISTERS_reg_67_16_inst : DFFR_X1 port map( D => n8476, CK => CLK, RN => 
                           n3012, Q => n10517, QN => n2239);
   REGISTERS_reg_67_15_inst : DFFR_X1 port map( D => n8477, CK => CLK, RN => 
                           n3012, Q => n10518, QN => n2240);
   REGISTERS_reg_67_14_inst : DFFR_X1 port map( D => n8478, CK => CLK, RN => 
                           n3012, Q => n10519, QN => n2241);
   REGISTERS_reg_67_13_inst : DFFR_X1 port map( D => n8479, CK => CLK, RN => 
                           n3012, Q => n10520, QN => n2242);
   REGISTERS_reg_67_12_inst : DFFR_X1 port map( D => n8480, CK => CLK, RN => 
                           n3012, Q => n10521, QN => n2243);
   REGISTERS_reg_67_11_inst : DFFR_X1 port map( D => n8481, CK => CLK, RN => 
                           n3011, Q => n10522, QN => n2244);
   REGISTERS_reg_67_10_inst : DFFR_X1 port map( D => n8482, CK => CLK, RN => 
                           n3011, Q => n10523, QN => n2245);
   REGISTERS_reg_67_9_inst : DFFR_X1 port map( D => n8483, CK => CLK, RN => 
                           n3011, Q => n10524, QN => n2246);
   REGISTERS_reg_67_8_inst : DFFR_X1 port map( D => n8484, CK => CLK, RN => 
                           n3011, Q => n10525, QN => n2247);
   REGISTERS_reg_67_7_inst : DFFR_X1 port map( D => n8485, CK => CLK, RN => 
                           n3011, Q => n10526, QN => n2248);
   REGISTERS_reg_67_6_inst : DFFR_X1 port map( D => n8486, CK => CLK, RN => 
                           n3011, Q => n10527, QN => n2249);
   REGISTERS_reg_67_5_inst : DFFR_X1 port map( D => n8487, CK => CLK, RN => 
                           n3011, Q => n10528, QN => n2250);
   REGISTERS_reg_67_4_inst : DFFR_X1 port map( D => n8488, CK => CLK, RN => 
                           n3011, Q => n10529, QN => n2251);
   REGISTERS_reg_67_3_inst : DFFR_X1 port map( D => n8489, CK => CLK, RN => 
                           n3011, Q => n10530, QN => n2252);
   REGISTERS_reg_67_2_inst : DFFR_X1 port map( D => n8490, CK => CLK, RN => 
                           n3011, Q => n10531, QN => n2253);
   REGISTERS_reg_67_1_inst : DFFR_X1 port map( D => n8491, CK => CLK, RN => 
                           n3011, Q => n10532, QN => n2254);
   REGISTERS_reg_67_0_inst : DFFR_X1 port map( D => n8492, CK => CLK, RN => 
                           n3011, Q => n10533, QN => n2255);
   REGISTERS_reg_68_31_inst : DFFR_X1 port map( D => n8493, CK => CLK, RN => 
                           n3010, Q => n10534, QN => n2256);
   REGISTERS_reg_68_30_inst : DFFR_X1 port map( D => n8494, CK => CLK, RN => 
                           n3010, Q => n10535, QN => n2257);
   REGISTERS_reg_68_29_inst : DFFR_X1 port map( D => n8495, CK => CLK, RN => 
                           n3010, Q => n10536, QN => n2258);
   REGISTERS_reg_68_28_inst : DFFR_X1 port map( D => n8496, CK => CLK, RN => 
                           n3010, Q => n10537, QN => n2259);
   REGISTERS_reg_68_27_inst : DFFR_X1 port map( D => n8497, CK => CLK, RN => 
                           n3010, Q => n10538, QN => n2260);
   REGISTERS_reg_68_26_inst : DFFR_X1 port map( D => n8498, CK => CLK, RN => 
                           n3010, Q => n10539, QN => n2261);
   REGISTERS_reg_68_25_inst : DFFR_X1 port map( D => n8499, CK => CLK, RN => 
                           n3010, Q => n10540, QN => n2262);
   REGISTERS_reg_68_24_inst : DFFR_X1 port map( D => n8500, CK => CLK, RN => 
                           n3010, Q => n10541, QN => n2263);
   REGISTERS_reg_68_23_inst : DFFR_X1 port map( D => n8501, CK => CLK, RN => 
                           n3010, Q => n10542, QN => n2264);
   REGISTERS_reg_68_22_inst : DFFR_X1 port map( D => n8502, CK => CLK, RN => 
                           n3010, Q => n10543, QN => n2265);
   REGISTERS_reg_68_21_inst : DFFR_X1 port map( D => n8503, CK => CLK, RN => 
                           n3010, Q => n10544, QN => n2266);
   REGISTERS_reg_68_20_inst : DFFR_X1 port map( D => n8504, CK => CLK, RN => 
                           n3010, Q => n10545, QN => n2267);
   REGISTERS_reg_68_19_inst : DFFR_X1 port map( D => n8505, CK => CLK, RN => 
                           n3009, Q => n10546, QN => n2268);
   REGISTERS_reg_68_18_inst : DFFR_X1 port map( D => n8506, CK => CLK, RN => 
                           n3009, Q => n10547, QN => n2269);
   REGISTERS_reg_68_17_inst : DFFR_X1 port map( D => n8507, CK => CLK, RN => 
                           n3009, Q => n10548, QN => n2270);
   REGISTERS_reg_68_16_inst : DFFR_X1 port map( D => n8508, CK => CLK, RN => 
                           n3009, Q => n10549, QN => n2271);
   REGISTERS_reg_68_15_inst : DFFR_X1 port map( D => n8509, CK => CLK, RN => 
                           n3009, Q => n10550, QN => n2272);
   REGISTERS_reg_68_14_inst : DFFR_X1 port map( D => n8510, CK => CLK, RN => 
                           n3009, Q => n10551, QN => n2273);
   REGISTERS_reg_68_13_inst : DFFR_X1 port map( D => n8511, CK => CLK, RN => 
                           n3009, Q => n10552, QN => n2274);
   REGISTERS_reg_68_12_inst : DFFR_X1 port map( D => n8512, CK => CLK, RN => 
                           n3009, Q => n10553, QN => n2275);
   REGISTERS_reg_68_11_inst : DFFR_X1 port map( D => n8513, CK => CLK, RN => 
                           n3009, Q => n10554, QN => n2276);
   REGISTERS_reg_68_10_inst : DFFR_X1 port map( D => n8514, CK => CLK, RN => 
                           n3009, Q => n10555, QN => n2277);
   REGISTERS_reg_68_9_inst : DFFR_X1 port map( D => n8515, CK => CLK, RN => 
                           n3009, Q => n10556, QN => n2278);
   REGISTERS_reg_68_8_inst : DFFR_X1 port map( D => n8516, CK => CLK, RN => 
                           n3009, Q => n10557, QN => n2279);
   REGISTERS_reg_68_7_inst : DFFR_X1 port map( D => n8517, CK => CLK, RN => 
                           n3008, Q => n10558, QN => n2280);
   REGISTERS_reg_68_6_inst : DFFR_X1 port map( D => n8518, CK => CLK, RN => 
                           n3008, Q => n10559, QN => n2281);
   REGISTERS_reg_68_5_inst : DFFR_X1 port map( D => n8519, CK => CLK, RN => 
                           n3008, Q => n10560, QN => n2282);
   REGISTERS_reg_68_4_inst : DFFR_X1 port map( D => n8520, CK => CLK, RN => 
                           n3008, Q => n10561, QN => n2283);
   REGISTERS_reg_68_3_inst : DFFR_X1 port map( D => n8521, CK => CLK, RN => 
                           n3008, Q => n10562, QN => n2284);
   REGISTERS_reg_68_2_inst : DFFR_X1 port map( D => n8522, CK => CLK, RN => 
                           n3008, Q => n10563, QN => n2285);
   REGISTERS_reg_68_1_inst : DFFR_X1 port map( D => n8523, CK => CLK, RN => 
                           n3008, Q => n10564, QN => n2286);
   REGISTERS_reg_68_0_inst : DFFR_X1 port map( D => n8524, CK => CLK, RN => 
                           n3008, Q => n10565, QN => n2287);
   REGISTERS_reg_69_31_inst : DFFR_X1 port map( D => n8525, CK => CLK, RN => 
                           n3008, Q => n10566, QN => n2288);
   REGISTERS_reg_69_30_inst : DFFR_X1 port map( D => n8526, CK => CLK, RN => 
                           n3008, Q => n10567, QN => n2289);
   REGISTERS_reg_69_29_inst : DFFR_X1 port map( D => n8527, CK => CLK, RN => 
                           n3008, Q => n10568, QN => n2290);
   REGISTERS_reg_69_28_inst : DFFR_X1 port map( D => n8528, CK => CLK, RN => 
                           n3008, Q => n10569, QN => n2291);
   REGISTERS_reg_69_27_inst : DFFR_X1 port map( D => n8529, CK => CLK, RN => 
                           n3007, Q => n10570, QN => n2292);
   REGISTERS_reg_69_26_inst : DFFR_X1 port map( D => n8530, CK => CLK, RN => 
                           n3007, Q => n10571, QN => n2293);
   REGISTERS_reg_69_25_inst : DFFR_X1 port map( D => n8531, CK => CLK, RN => 
                           n3007, Q => n10572, QN => n2294);
   REGISTERS_reg_69_24_inst : DFFR_X1 port map( D => n8532, CK => CLK, RN => 
                           n3007, Q => n10573, QN => n2295);
   REGISTERS_reg_69_23_inst : DFFR_X1 port map( D => n8533, CK => CLK, RN => 
                           n3007, Q => n10574, QN => n2296);
   REGISTERS_reg_69_22_inst : DFFR_X1 port map( D => n8534, CK => CLK, RN => 
                           n3007, Q => n10575, QN => n2297);
   REGISTERS_reg_69_21_inst : DFFR_X1 port map( D => n8535, CK => CLK, RN => 
                           n3007, Q => n10576, QN => n2298);
   REGISTERS_reg_69_20_inst : DFFR_X1 port map( D => n8536, CK => CLK, RN => 
                           n3007, Q => n10577, QN => n2299);
   REGISTERS_reg_69_19_inst : DFFR_X1 port map( D => n8537, CK => CLK, RN => 
                           n3007, Q => n10578, QN => n2300);
   REGISTERS_reg_69_18_inst : DFFR_X1 port map( D => n8538, CK => CLK, RN => 
                           n3007, Q => n10579, QN => n2301);
   REGISTERS_reg_69_17_inst : DFFR_X1 port map( D => n8539, CK => CLK, RN => 
                           n3007, Q => n10580, QN => n2302);
   REGISTERS_reg_69_16_inst : DFFR_X1 port map( D => n8540, CK => CLK, RN => 
                           n3007, Q => n10581, QN => n2303);
   REGISTERS_reg_69_15_inst : DFFR_X1 port map( D => n8541, CK => CLK, RN => 
                           n3006, Q => n10582, QN => n2304);
   REGISTERS_reg_69_14_inst : DFFR_X1 port map( D => n8542, CK => CLK, RN => 
                           n3006, Q => n10583, QN => n2305);
   REGISTERS_reg_69_13_inst : DFFR_X1 port map( D => n8543, CK => CLK, RN => 
                           n3006, Q => n10584, QN => n2306);
   REGISTERS_reg_69_12_inst : DFFR_X1 port map( D => n8544, CK => CLK, RN => 
                           n3006, Q => n10585, QN => n2307);
   REGISTERS_reg_69_11_inst : DFFR_X1 port map( D => n8545, CK => CLK, RN => 
                           n3006, Q => n10586, QN => n2308);
   REGISTERS_reg_69_10_inst : DFFR_X1 port map( D => n8546, CK => CLK, RN => 
                           n3006, Q => n10587, QN => n2309);
   REGISTERS_reg_69_9_inst : DFFR_X1 port map( D => n8547, CK => CLK, RN => 
                           n3006, Q => n10588, QN => n2310);
   REGISTERS_reg_69_8_inst : DFFR_X1 port map( D => n8548, CK => CLK, RN => 
                           n3006, Q => n10589, QN => n2311);
   REGISTERS_reg_69_7_inst : DFFR_X1 port map( D => n8549, CK => CLK, RN => 
                           n3006, Q => n10590, QN => n2312);
   REGISTERS_reg_69_6_inst : DFFR_X1 port map( D => n8550, CK => CLK, RN => 
                           n3006, Q => n10591, QN => n2313);
   REGISTERS_reg_69_5_inst : DFFR_X1 port map( D => n8551, CK => CLK, RN => 
                           n3006, Q => n10592, QN => n2314);
   REGISTERS_reg_69_4_inst : DFFR_X1 port map( D => n8552, CK => CLK, RN => 
                           n3006, Q => n10593, QN => n2315);
   REGISTERS_reg_69_3_inst : DFFR_X1 port map( D => n8553, CK => CLK, RN => 
                           n3005, Q => n10594, QN => n2316);
   REGISTERS_reg_69_2_inst : DFFR_X1 port map( D => n8554, CK => CLK, RN => 
                           n3005, Q => n10595, QN => n2317);
   REGISTERS_reg_69_1_inst : DFFR_X1 port map( D => n8555, CK => CLK, RN => 
                           n3005, Q => n10596, QN => n2318);
   REGISTERS_reg_69_0_inst : DFFR_X1 port map( D => n8556, CK => CLK, RN => 
                           n3005, Q => n10597, QN => n2319);
   REGISTERS_reg_70_31_inst : DFFR_X1 port map( D => n8557, CK => CLK, RN => 
                           n3005, Q => n10598, QN => n2320);
   REGISTERS_reg_70_30_inst : DFFR_X1 port map( D => n8558, CK => CLK, RN => 
                           n3005, Q => n10599, QN => n2321);
   REGISTERS_reg_70_29_inst : DFFR_X1 port map( D => n8559_port, CK => CLK, RN 
                           => n3005, Q => n10600, QN => n2322);
   REGISTERS_reg_70_28_inst : DFFR_X1 port map( D => n8560, CK => CLK, RN => 
                           n3005, Q => n10601, QN => n2323);
   REGISTERS_reg_70_27_inst : DFFR_X1 port map( D => n8561_port, CK => CLK, RN 
                           => n3005, Q => n10602, QN => n2324);
   REGISTERS_reg_70_26_inst : DFFR_X1 port map( D => n8562_port, CK => CLK, RN 
                           => n3005, Q => n10603, QN => n2325);
   REGISTERS_reg_70_25_inst : DFFR_X1 port map( D => n8563_port, CK => CLK, RN 
                           => n3005, Q => n10604, QN => n2326);
   REGISTERS_reg_70_24_inst : DFFR_X1 port map( D => n8564_port, CK => CLK, RN 
                           => n3005, Q => n10605, QN => n2327);
   REGISTERS_reg_70_23_inst : DFFR_X1 port map( D => n8565_port, CK => CLK, RN 
                           => n3004, Q => n10606, QN => n2328);
   REGISTERS_reg_70_22_inst : DFFR_X1 port map( D => n8566_port, CK => CLK, RN 
                           => n3004, Q => n10607, QN => n2329);
   REGISTERS_reg_70_21_inst : DFFR_X1 port map( D => n8567_port, CK => CLK, RN 
                           => n3004, Q => n10608, QN => n2330);
   REGISTERS_reg_70_20_inst : DFFR_X1 port map( D => n8568, CK => CLK, RN => 
                           n3004, Q => n10609, QN => n2331);
   REGISTERS_reg_70_19_inst : DFFR_X1 port map( D => n8569, CK => CLK, RN => 
                           n3004, Q => n10610, QN => n2332);
   REGISTERS_reg_70_18_inst : DFFR_X1 port map( D => n8570, CK => CLK, RN => 
                           n3004, Q => n10611, QN => n2333);
   REGISTERS_reg_70_17_inst : DFFR_X1 port map( D => n8571_port, CK => CLK, RN 
                           => n3004, Q => n10612, QN => n2334);
   REGISTERS_reg_70_16_inst : DFFR_X1 port map( D => n8572_port, CK => CLK, RN 
                           => n3004, Q => n10613, QN => n2335);
   REGISTERS_reg_70_15_inst : DFFR_X1 port map( D => n8573_port, CK => CLK, RN 
                           => n3004, Q => n10614, QN => n2336);
   REGISTERS_reg_70_14_inst : DFFR_X1 port map( D => n8574_port, CK => CLK, RN 
                           => n3004, Q => n10615, QN => n2337);
   REGISTERS_reg_70_13_inst : DFFR_X1 port map( D => n8575, CK => CLK, RN => 
                           n3004, Q => n10616, QN => n2338);
   REGISTERS_reg_70_12_inst : DFFR_X1 port map( D => n8576, CK => CLK, RN => 
                           n3004, Q => n10617, QN => n2339);
   REGISTERS_reg_70_11_inst : DFFR_X1 port map( D => n8577, CK => CLK, RN => 
                           n3003, Q => n10618, QN => n2340);
   REGISTERS_reg_70_10_inst : DFFR_X1 port map( D => n8578, CK => CLK, RN => 
                           n3003, Q => n10619, QN => n2341);
   REGISTERS_reg_70_9_inst : DFFR_X1 port map( D => n8579, CK => CLK, RN => 
                           n3003, Q => n10620, QN => n2342);
   REGISTERS_reg_70_8_inst : DFFR_X1 port map( D => n8580, CK => CLK, RN => 
                           n3003, Q => n10621, QN => n2343);
   REGISTERS_reg_70_7_inst : DFFR_X1 port map( D => n8581, CK => CLK, RN => 
                           n3003, Q => n10622, QN => n2344);
   REGISTERS_reg_70_6_inst : DFFR_X1 port map( D => n8582, CK => CLK, RN => 
                           n3003, Q => n10623, QN => n2345);
   REGISTERS_reg_70_5_inst : DFFR_X1 port map( D => n8583, CK => CLK, RN => 
                           n3003, Q => n10624, QN => n2346);
   REGISTERS_reg_70_4_inst : DFFR_X1 port map( D => n8584, CK => CLK, RN => 
                           n3003, Q => n10625, QN => n2347);
   REGISTERS_reg_70_3_inst : DFFR_X1 port map( D => n8585, CK => CLK, RN => 
                           n3003, Q => n10626, QN => n2348);
   REGISTERS_reg_70_2_inst : DFFR_X1 port map( D => n8586, CK => CLK, RN => 
                           n3003, Q => n10627, QN => n2349);
   REGISTERS_reg_70_1_inst : DFFR_X1 port map( D => n8587, CK => CLK, RN => 
                           n3003, Q => n10628, QN => n2350);
   REGISTERS_reg_70_0_inst : DFFR_X1 port map( D => n8588, CK => CLK, RN => 
                           n3003, Q => n10629, QN => n2351);
   REGISTERS_reg_71_31_inst : DFFR_X1 port map( D => n8589, CK => CLK, RN => 
                           n3002, Q => n10630, QN => n2352);
   REGISTERS_reg_71_30_inst : DFFR_X1 port map( D => n8590, CK => CLK, RN => 
                           n3002, Q => n10631, QN => n2353);
   REGISTERS_reg_71_29_inst : DFFR_X1 port map( D => n8591, CK => CLK, RN => 
                           n3002, Q => n10632, QN => n2354);
   REGISTERS_reg_71_28_inst : DFFR_X1 port map( D => n8592, CK => CLK, RN => 
                           n3002, Q => n10633, QN => n2355);
   REGISTERS_reg_71_27_inst : DFFR_X1 port map( D => n8593, CK => CLK, RN => 
                           n3002, Q => n10634, QN => n2356);
   REGISTERS_reg_71_26_inst : DFFR_X1 port map( D => n8594, CK => CLK, RN => 
                           n3002, Q => n10635, QN => n2357);
   REGISTERS_reg_71_25_inst : DFFR_X1 port map( D => n8595, CK => CLK, RN => 
                           n3002, Q => n10636, QN => n2358);
   REGISTERS_reg_71_24_inst : DFFR_X1 port map( D => n8596, CK => CLK, RN => 
                           n3002, Q => n10637, QN => n2359);
   REGISTERS_reg_71_23_inst : DFFR_X1 port map( D => n8597, CK => CLK, RN => 
                           n3002, Q => n10638, QN => n2360);
   REGISTERS_reg_71_22_inst : DFFR_X1 port map( D => n8598, CK => CLK, RN => 
                           n3002, Q => n10639, QN => n2361);
   REGISTERS_reg_71_21_inst : DFFR_X1 port map( D => n8599, CK => CLK, RN => 
                           n3002, Q => n10640, QN => n2362);
   REGISTERS_reg_71_20_inst : DFFR_X1 port map( D => n8600, CK => CLK, RN => 
                           n3002, Q => n10641, QN => n2363);
   REGISTERS_reg_71_19_inst : DFFR_X1 port map( D => n8601, CK => CLK, RN => 
                           n3001, Q => n10642, QN => n2364);
   REGISTERS_reg_71_18_inst : DFFR_X1 port map( D => n8602, CK => CLK, RN => 
                           n3001, Q => n10643, QN => n2365);
   REGISTERS_reg_71_17_inst : DFFR_X1 port map( D => n8603, CK => CLK, RN => 
                           n3001, Q => n10644, QN => n2366);
   REGISTERS_reg_71_16_inst : DFFR_X1 port map( D => n8604, CK => CLK, RN => 
                           n3001, Q => n10645, QN => n2367);
   REGISTERS_reg_71_15_inst : DFFR_X1 port map( D => n8605, CK => CLK, RN => 
                           n3001, Q => n10646, QN => n2368);
   REGISTERS_reg_71_14_inst : DFFR_X1 port map( D => n8606, CK => CLK, RN => 
                           n3001, Q => n10647, QN => n2369);
   REGISTERS_reg_71_13_inst : DFFR_X1 port map( D => n8607, CK => CLK, RN => 
                           n3001, Q => n10648, QN => n2370);
   REGISTERS_reg_71_12_inst : DFFR_X1 port map( D => n8608, CK => CLK, RN => 
                           n3001, Q => n10649, QN => n2371);
   REGISTERS_reg_71_11_inst : DFFR_X1 port map( D => n8609, CK => CLK, RN => 
                           n3001, Q => n10650, QN => n2372);
   REGISTERS_reg_71_10_inst : DFFR_X1 port map( D => n8610, CK => CLK, RN => 
                           n3001, Q => n10651, QN => n2373);
   REGISTERS_reg_71_9_inst : DFFR_X1 port map( D => n8611, CK => CLK, RN => 
                           n3001, Q => n10652, QN => n2374);
   REGISTERS_reg_71_8_inst : DFFR_X1 port map( D => n8612, CK => CLK, RN => 
                           n3001, Q => n10653, QN => n2375);
   REGISTERS_reg_71_7_inst : DFFR_X1 port map( D => n8613, CK => CLK, RN => 
                           n3000, Q => n10654, QN => n2376);
   REGISTERS_reg_71_6_inst : DFFR_X1 port map( D => n8614, CK => CLK, RN => 
                           n3000, Q => n10655, QN => n2377);
   REGISTERS_reg_71_5_inst : DFFR_X1 port map( D => n8615, CK => CLK, RN => 
                           n3000, Q => n10656, QN => n2378);
   REGISTERS_reg_71_4_inst : DFFR_X1 port map( D => n8616, CK => CLK, RN => 
                           n3000, Q => n10657, QN => n2379);
   REGISTERS_reg_71_3_inst : DFFR_X1 port map( D => n8617, CK => CLK, RN => 
                           n3000, Q => n10658, QN => n2380);
   REGISTERS_reg_71_2_inst : DFFR_X1 port map( D => n8618, CK => CLK, RN => 
                           n3000, Q => n10659, QN => n2381);
   REGISTERS_reg_71_1_inst : DFFR_X1 port map( D => n8619, CK => CLK, RN => 
                           n3000, Q => n10660, QN => n2382);
   REGISTERS_reg_71_0_inst : DFFR_X1 port map( D => n8620, CK => CLK, RN => 
                           n3000, Q => n10661, QN => n2383);
   REGISTERS_reg_72_31_inst : DFFR_X1 port map( D => n8621, CK => CLK, RN => 
                           n3000, Q => n10662, QN => n2384);
   REGISTERS_reg_72_30_inst : DFFR_X1 port map( D => n8622, CK => CLK, RN => 
                           n3000, Q => n10663, QN => n2385);
   REGISTERS_reg_72_29_inst : DFFR_X1 port map( D => n8623, CK => CLK, RN => 
                           n3000, Q => n10664, QN => n2386);
   REGISTERS_reg_72_28_inst : DFFR_X1 port map( D => n8624, CK => CLK, RN => 
                           n3000, Q => n10665, QN => n2387);
   REGISTERS_reg_72_27_inst : DFFR_X1 port map( D => n8625, CK => CLK, RN => 
                           n2999, Q => n10666, QN => n2388);
   REGISTERS_reg_72_26_inst : DFFR_X1 port map( D => n8626, CK => CLK, RN => 
                           n2999, Q => n10667, QN => n2389);
   REGISTERS_reg_72_25_inst : DFFR_X1 port map( D => n8627, CK => CLK, RN => 
                           n2999, Q => n10668, QN => n2390);
   REGISTERS_reg_72_24_inst : DFFR_X1 port map( D => n8628, CK => CLK, RN => 
                           n2999, Q => n10669, QN => n2391);
   REGISTERS_reg_72_23_inst : DFFR_X1 port map( D => n8629, CK => CLK, RN => 
                           n2999, Q => n10670, QN => n2392);
   REGISTERS_reg_72_22_inst : DFFR_X1 port map( D => n8630, CK => CLK, RN => 
                           n2999, Q => n10671, QN => n2393);
   REGISTERS_reg_72_21_inst : DFFR_X1 port map( D => n8631, CK => CLK, RN => 
                           n2999, Q => n10672, QN => n2394);
   REGISTERS_reg_72_20_inst : DFFR_X1 port map( D => n8632, CK => CLK, RN => 
                           n2999, Q => n10673, QN => n2395);
   REGISTERS_reg_72_19_inst : DFFR_X1 port map( D => n8633, CK => CLK, RN => 
                           n2999, Q => n10674, QN => n2396);
   REGISTERS_reg_72_18_inst : DFFR_X1 port map( D => n8634, CK => CLK, RN => 
                           n2999, Q => n10675, QN => n2397);
   REGISTERS_reg_72_17_inst : DFFR_X1 port map( D => n8635, CK => CLK, RN => 
                           n2999, Q => n10676, QN => n2398);
   REGISTERS_reg_72_16_inst : DFFR_X1 port map( D => n8636, CK => CLK, RN => 
                           n2999, Q => n10677, QN => n2399);
   REGISTERS_reg_72_15_inst : DFFR_X1 port map( D => n8637, CK => CLK, RN => 
                           n2998, Q => n10678, QN => n2400);
   REGISTERS_reg_72_14_inst : DFFR_X1 port map( D => n8638, CK => CLK, RN => 
                           n2998, Q => n10679, QN => n2401);
   REGISTERS_reg_72_13_inst : DFFR_X1 port map( D => n8639, CK => CLK, RN => 
                           n2998, Q => n10680, QN => n2402);
   REGISTERS_reg_72_12_inst : DFFR_X1 port map( D => n8640, CK => CLK, RN => 
                           n2998, Q => n10681, QN => n2403);
   REGISTERS_reg_72_11_inst : DFFR_X1 port map( D => n8641, CK => CLK, RN => 
                           n2998, Q => n10682, QN => n2404);
   REGISTERS_reg_72_10_inst : DFFR_X1 port map( D => n8642, CK => CLK, RN => 
                           n2998, Q => n10683, QN => n2405);
   REGISTERS_reg_72_9_inst : DFFR_X1 port map( D => n8643, CK => CLK, RN => 
                           n2998, Q => n10684, QN => n2406);
   REGISTERS_reg_72_8_inst : DFFR_X1 port map( D => n8644, CK => CLK, RN => 
                           n2998, Q => n10685, QN => n2407);
   REGISTERS_reg_72_7_inst : DFFR_X1 port map( D => n8645, CK => CLK, RN => 
                           n2998, Q => n10686, QN => n2408);
   REGISTERS_reg_72_6_inst : DFFR_X1 port map( D => n8646, CK => CLK, RN => 
                           n2998, Q => n10687, QN => n2409);
   REGISTERS_reg_72_5_inst : DFFR_X1 port map( D => n8647, CK => CLK, RN => 
                           n2998, Q => n10688, QN => n2410);
   REGISTERS_reg_72_4_inst : DFFR_X1 port map( D => n8648, CK => CLK, RN => 
                           n2998, Q => n10689, QN => n2411);
   REGISTERS_reg_72_3_inst : DFFR_X1 port map( D => n8649, CK => CLK, RN => 
                           n2997, Q => n10690, QN => n2412);
   REGISTERS_reg_72_2_inst : DFFR_X1 port map( D => n8650, CK => CLK, RN => 
                           n2997, Q => n10691, QN => n2413);
   REGISTERS_reg_72_1_inst : DFFR_X1 port map( D => n8651, CK => CLK, RN => 
                           n2997, Q => n10692, QN => n2414);
   REGISTERS_reg_72_0_inst : DFFR_X1 port map( D => n8652, CK => CLK, RN => 
                           n2997, Q => n10693, QN => n2415);
   REGISTERS_reg_73_31_inst : DFFR_X1 port map( D => n8653, CK => CLK, RN => 
                           n2997, Q => n10694, QN => n2416);
   REGISTERS_reg_73_30_inst : DFFR_X1 port map( D => n8654, CK => CLK, RN => 
                           n2997, Q => n10695, QN => n2417);
   REGISTERS_reg_73_29_inst : DFFR_X1 port map( D => n8655, CK => CLK, RN => 
                           n2997, Q => n10696, QN => n2418);
   REGISTERS_reg_73_28_inst : DFFR_X1 port map( D => n8656, CK => CLK, RN => 
                           n2997, Q => n10697, QN => n2419);
   REGISTERS_reg_73_27_inst : DFFR_X1 port map( D => n8657, CK => CLK, RN => 
                           n2997, Q => n10698, QN => n2420);
   REGISTERS_reg_73_26_inst : DFFR_X1 port map( D => n8658, CK => CLK, RN => 
                           n2997, Q => n10699, QN => n2421);
   REGISTERS_reg_73_25_inst : DFFR_X1 port map( D => n8659, CK => CLK, RN => 
                           n2997, Q => n10700, QN => n2422);
   REGISTERS_reg_73_24_inst : DFFR_X1 port map( D => n8660, CK => CLK, RN => 
                           n2997, Q => n10701, QN => n2423);
   REGISTERS_reg_73_23_inst : DFFR_X1 port map( D => n8661, CK => CLK, RN => 
                           n2995, Q => n10702, QN => n2424);
   REGISTERS_reg_73_22_inst : DFFR_X1 port map( D => n8662, CK => CLK, RN => 
                           n2995, Q => n10703, QN => n2425);
   REGISTERS_reg_73_21_inst : DFFR_X1 port map( D => n8663, CK => CLK, RN => 
                           n2995, Q => n10704, QN => n2426);
   REGISTERS_reg_73_20_inst : DFFR_X1 port map( D => n8664, CK => CLK, RN => 
                           n2995, Q => n10705, QN => n2427);
   REGISTERS_reg_73_19_inst : DFFR_X1 port map( D => n8665, CK => CLK, RN => 
                           n2995, Q => n10706, QN => n2428);
   REGISTERS_reg_73_18_inst : DFFR_X1 port map( D => n8666, CK => CLK, RN => 
                           n2995, Q => n10707, QN => n2429);
   REGISTERS_reg_73_17_inst : DFFR_X1 port map( D => n8667, CK => CLK, RN => 
                           n2995, Q => n10708, QN => n2430);
   REGISTERS_reg_73_16_inst : DFFR_X1 port map( D => n8668, CK => CLK, RN => 
                           n2995, Q => n10709, QN => n2431);
   REGISTERS_reg_73_15_inst : DFFR_X1 port map( D => n8669, CK => CLK, RN => 
                           n2995, Q => n10710, QN => n2432);
   REGISTERS_reg_73_14_inst : DFFR_X1 port map( D => n8670, CK => CLK, RN => 
                           n2995, Q => n10711, QN => n2433);
   REGISTERS_reg_73_13_inst : DFFR_X1 port map( D => n8671, CK => CLK, RN => 
                           n2995, Q => n10712, QN => n2434);
   REGISTERS_reg_73_12_inst : DFFR_X1 port map( D => n8672, CK => CLK, RN => 
                           n2995, Q => n10713, QN => n2435);
   REGISTERS_reg_73_11_inst : DFFR_X1 port map( D => n8673, CK => CLK, RN => 
                           n2994, Q => n10714, QN => n2436);
   REGISTERS_reg_73_10_inst : DFFR_X1 port map( D => n8674, CK => CLK, RN => 
                           n2994, Q => n10715, QN => n2437);
   REGISTERS_reg_73_9_inst : DFFR_X1 port map( D => n8675, CK => CLK, RN => 
                           n2994, Q => n10716, QN => n2438);
   REGISTERS_reg_73_8_inst : DFFR_X1 port map( D => n8676, CK => CLK, RN => 
                           n2994, Q => n10717, QN => n2439);
   REGISTERS_reg_73_7_inst : DFFR_X1 port map( D => n8677, CK => CLK, RN => 
                           n2994, Q => n10718, QN => n2440);
   REGISTERS_reg_73_6_inst : DFFR_X1 port map( D => n8678, CK => CLK, RN => 
                           n2994, Q => n10719, QN => n2441);
   REGISTERS_reg_73_5_inst : DFFR_X1 port map( D => n8679, CK => CLK, RN => 
                           n2994, Q => n10720, QN => n2442);
   REGISTERS_reg_73_4_inst : DFFR_X1 port map( D => n8680, CK => CLK, RN => 
                           n2994, Q => n10721, QN => n2443);
   REGISTERS_reg_73_3_inst : DFFR_X1 port map( D => n8681, CK => CLK, RN => 
                           n2994, Q => n10722, QN => n2444);
   REGISTERS_reg_73_2_inst : DFFR_X1 port map( D => n8682, CK => CLK, RN => 
                           n2994, Q => n10723, QN => n2445);
   REGISTERS_reg_73_1_inst : DFFR_X1 port map( D => n8683, CK => CLK, RN => 
                           n2994, Q => n10724, QN => n2446);
   REGISTERS_reg_73_0_inst : DFFR_X1 port map( D => n8684, CK => CLK, RN => 
                           n2994, Q => n10725, QN => n2447);
   REGISTERS_reg_74_31_inst : DFFR_X1 port map( D => n8685, CK => CLK, RN => 
                           n2993, Q => n10726, QN => n2448);
   REGISTERS_reg_74_30_inst : DFFR_X1 port map( D => n8686, CK => CLK, RN => 
                           n2993, Q => n10727, QN => n2449);
   REGISTERS_reg_74_29_inst : DFFR_X1 port map( D => n8687, CK => CLK, RN => 
                           n2993, Q => n10728, QN => n2450);
   REGISTERS_reg_74_28_inst : DFFR_X1 port map( D => n8688, CK => CLK, RN => 
                           n2993, Q => n10729, QN => n2451);
   REGISTERS_reg_74_27_inst : DFFR_X1 port map( D => n8689, CK => CLK, RN => 
                           n2993, Q => n10730, QN => n2452);
   REGISTERS_reg_74_26_inst : DFFR_X1 port map( D => n8690, CK => CLK, RN => 
                           n2993, Q => n10731, QN => n2453);
   REGISTERS_reg_74_25_inst : DFFR_X1 port map( D => n8691, CK => CLK, RN => 
                           n2993, Q => n10732, QN => n2454);
   REGISTERS_reg_74_24_inst : DFFR_X1 port map( D => n8692, CK => CLK, RN => 
                           n2993, Q => n10733, QN => n2455);
   REGISTERS_reg_74_23_inst : DFFR_X1 port map( D => n8693, CK => CLK, RN => 
                           n2993, Q => n10734, QN => n2456);
   REGISTERS_reg_74_22_inst : DFFR_X1 port map( D => n8694, CK => CLK, RN => 
                           n2993, Q => n10735, QN => n2457);
   REGISTERS_reg_74_21_inst : DFFR_X1 port map( D => n8695, CK => CLK, RN => 
                           n2993, Q => n10736, QN => n2458);
   REGISTERS_reg_74_20_inst : DFFR_X1 port map( D => n8696, CK => CLK, RN => 
                           n2993, Q => n10737, QN => n2459);
   REGISTERS_reg_74_19_inst : DFFR_X1 port map( D => n8697, CK => CLK, RN => 
                           n2992, Q => n10738, QN => n2460);
   REGISTERS_reg_74_18_inst : DFFR_X1 port map( D => n8698, CK => CLK, RN => 
                           n2992, Q => n10739, QN => n2461);
   REGISTERS_reg_74_17_inst : DFFR_X1 port map( D => n8699, CK => CLK, RN => 
                           n2992, Q => n10740, QN => n2462);
   REGISTERS_reg_74_16_inst : DFFR_X1 port map( D => n8700, CK => CLK, RN => 
                           n2992, Q => n10741, QN => n2463);
   REGISTERS_reg_74_15_inst : DFFR_X1 port map( D => n8701, CK => CLK, RN => 
                           n2992, Q => n10742, QN => n2464);
   REGISTERS_reg_74_14_inst : DFFR_X1 port map( D => n8702_port, CK => CLK, RN 
                           => n2992, Q => n10743, QN => n2465);
   REGISTERS_reg_74_13_inst : DFFR_X1 port map( D => n8703_port, CK => CLK, RN 
                           => n2992, Q => n10744, QN => n2466);
   REGISTERS_reg_74_12_inst : DFFR_X1 port map( D => n8704_port, CK => CLK, RN 
                           => n2992, Q => n10745, QN => n2467);
   REGISTERS_reg_74_11_inst : DFFR_X1 port map( D => n8705_port, CK => CLK, RN 
                           => n2992, Q => n10746, QN => n2468);
   REGISTERS_reg_74_10_inst : DFFR_X1 port map( D => n8706_port, CK => CLK, RN 
                           => n2992, Q => n10747, QN => n2469);
   REGISTERS_reg_74_9_inst : DFFR_X1 port map( D => n8707_port, CK => CLK, RN 
                           => n2992, Q => n10748, QN => n2470);
   REGISTERS_reg_74_8_inst : DFFR_X1 port map( D => n8708_port, CK => CLK, RN 
                           => n2992, Q => n10749, QN => n2471);
   REGISTERS_reg_74_7_inst : DFFR_X1 port map( D => n8709_port, CK => CLK, RN 
                           => n2991, Q => n10750, QN => n2472);
   REGISTERS_reg_74_6_inst : DFFR_X1 port map( D => n8710_port, CK => CLK, RN 
                           => n2991, Q => n10751, QN => n2473);
   REGISTERS_reg_74_5_inst : DFFR_X1 port map( D => n8711_port, CK => CLK, RN 
                           => n2991, Q => n10752, QN => n2474);
   REGISTERS_reg_74_4_inst : DFFR_X1 port map( D => n8712_port, CK => CLK, RN 
                           => n2991, Q => n10753, QN => n2475);
   REGISTERS_reg_74_3_inst : DFFR_X1 port map( D => n8713_port, CK => CLK, RN 
                           => n2991, Q => n10754, QN => n2476);
   REGISTERS_reg_74_2_inst : DFFR_X1 port map( D => n8714_port, CK => CLK, RN 
                           => n2991, Q => n10755, QN => n2477);
   REGISTERS_reg_74_1_inst : DFFR_X1 port map( D => n8715_port, CK => CLK, RN 
                           => n2991, Q => n10756, QN => n2478);
   REGISTERS_reg_74_0_inst : DFFR_X1 port map( D => n8716_port, CK => CLK, RN 
                           => n2991, Q => n10757, QN => n2479);
   REGISTERS_reg_75_31_inst : DFFR_X1 port map( D => n8717_port, CK => CLK, RN 
                           => n2991, Q => n10758, QN => n2480);
   REGISTERS_reg_75_30_inst : DFFR_X1 port map( D => n8718_port, CK => CLK, RN 
                           => n2991, Q => n10759, QN => n2481);
   REGISTERS_reg_75_29_inst : DFFR_X1 port map( D => n8719_port, CK => CLK, RN 
                           => n2991, Q => n10760, QN => n2482);
   REGISTERS_reg_75_28_inst : DFFR_X1 port map( D => n8720_port, CK => CLK, RN 
                           => n2991, Q => n10761, QN => n2483);
   REGISTERS_reg_75_27_inst : DFFR_X1 port map( D => n8721_port, CK => CLK, RN 
                           => n2990, Q => n10762, QN => n2484);
   REGISTERS_reg_75_26_inst : DFFR_X1 port map( D => n8722_port, CK => CLK, RN 
                           => n2990, Q => n10763, QN => n2485);
   REGISTERS_reg_75_25_inst : DFFR_X1 port map( D => n8723_port, CK => CLK, RN 
                           => n2990, Q => n10764, QN => n2486);
   REGISTERS_reg_75_24_inst : DFFR_X1 port map( D => n8724_port, CK => CLK, RN 
                           => n2990, Q => n10765, QN => n2487);
   REGISTERS_reg_75_23_inst : DFFR_X1 port map( D => n8725_port, CK => CLK, RN 
                           => n2990, Q => n10766, QN => n2488);
   REGISTERS_reg_75_22_inst : DFFR_X1 port map( D => n8726_port, CK => CLK, RN 
                           => n2990, Q => n10767, QN => n2489);
   REGISTERS_reg_75_21_inst : DFFR_X1 port map( D => n8727_port, CK => CLK, RN 
                           => n2990, Q => n10768, QN => n2490);
   REGISTERS_reg_75_20_inst : DFFR_X1 port map( D => n8728_port, CK => CLK, RN 
                           => n2990, Q => n10769, QN => n2491);
   REGISTERS_reg_75_19_inst : DFFR_X1 port map( D => n8729_port, CK => CLK, RN 
                           => n2990, Q => n10770, QN => n2492);
   REGISTERS_reg_75_18_inst : DFFR_X1 port map( D => n8730_port, CK => CLK, RN 
                           => n2990, Q => n10771, QN => n2493);
   REGISTERS_reg_75_17_inst : DFFR_X1 port map( D => n8731_port, CK => CLK, RN 
                           => n2990, Q => n10772, QN => n2494);
   REGISTERS_reg_75_16_inst : DFFR_X1 port map( D => n8732_port, CK => CLK, RN 
                           => n2990, Q => n10773, QN => n2495);
   REGISTERS_reg_75_15_inst : DFFR_X1 port map( D => n8733_port, CK => CLK, RN 
                           => n2989, Q => n10774, QN => n2496);
   REGISTERS_reg_75_14_inst : DFFR_X1 port map( D => n8734_port, CK => CLK, RN 
                           => n2989, Q => n10775, QN => n2497);
   REGISTERS_reg_75_13_inst : DFFR_X1 port map( D => n8735_port, CK => CLK, RN 
                           => n2989, Q => n10776, QN => n2498);
   REGISTERS_reg_75_12_inst : DFFR_X1 port map( D => n8736_port, CK => CLK, RN 
                           => n2989, Q => n10777, QN => n2499);
   REGISTERS_reg_75_11_inst : DFFR_X1 port map( D => n8737_port, CK => CLK, RN 
                           => n2989, Q => n10778, QN => n2500);
   REGISTERS_reg_75_10_inst : DFFR_X1 port map( D => n8738_port, CK => CLK, RN 
                           => n2989, Q => n10779, QN => n2501);
   REGISTERS_reg_75_9_inst : DFFR_X1 port map( D => n8739_port, CK => CLK, RN 
                           => n2989, Q => n10780, QN => n2502);
   REGISTERS_reg_75_8_inst : DFFR_X1 port map( D => n8740_port, CK => CLK, RN 
                           => n2989, Q => n10781, QN => n2503);
   REGISTERS_reg_75_7_inst : DFFR_X1 port map( D => n8741_port, CK => CLK, RN 
                           => n2989, Q => n10782, QN => n2504);
   REGISTERS_reg_75_6_inst : DFFR_X1 port map( D => n8742_port, CK => CLK, RN 
                           => n2989, Q => n10783, QN => n2505);
   REGISTERS_reg_75_5_inst : DFFR_X1 port map( D => n8743_port, CK => CLK, RN 
                           => n2989, Q => n10784, QN => n2506);
   REGISTERS_reg_75_4_inst : DFFR_X1 port map( D => n8744_port, CK => CLK, RN 
                           => n2989, Q => n10785, QN => n2507);
   REGISTERS_reg_75_3_inst : DFFR_X1 port map( D => n8745_port, CK => CLK, RN 
                           => n2988, Q => n10786, QN => n2508);
   REGISTERS_reg_75_2_inst : DFFR_X1 port map( D => n8746_port, CK => CLK, RN 
                           => n2988, Q => n10787, QN => n2509);
   REGISTERS_reg_75_1_inst : DFFR_X1 port map( D => n8747_port, CK => CLK, RN 
                           => n2988, Q => n10788, QN => n2510);
   REGISTERS_reg_75_0_inst : DFFR_X1 port map( D => n8748_port, CK => CLK, RN 
                           => n2988, Q => n10789, QN => n2511);
   REGISTERS_reg_76_31_inst : DFFR_X1 port map( D => n8749_port, CK => CLK, RN 
                           => n2988, Q => n10790, QN => n2512);
   REGISTERS_reg_76_30_inst : DFFR_X1 port map( D => n8750_port, CK => CLK, RN 
                           => n2988, Q => n10791, QN => n2513);
   REGISTERS_reg_76_29_inst : DFFR_X1 port map( D => n8751_port, CK => CLK, RN 
                           => n2988, Q => n10792, QN => n2514);
   REGISTERS_reg_76_28_inst : DFFR_X1 port map( D => n8752_port, CK => CLK, RN 
                           => n2988, Q => n10793, QN => n2515);
   REGISTERS_reg_76_27_inst : DFFR_X1 port map( D => n8753_port, CK => CLK, RN 
                           => n2988, Q => n10794, QN => n2516);
   REGISTERS_reg_76_26_inst : DFFR_X1 port map( D => n8754_port, CK => CLK, RN 
                           => n2988, Q => n10795, QN => n2517);
   REGISTERS_reg_76_25_inst : DFFR_X1 port map( D => n8755_port, CK => CLK, RN 
                           => n2988, Q => n10796, QN => n2518);
   REGISTERS_reg_76_24_inst : DFFR_X1 port map( D => n8756_port, CK => CLK, RN 
                           => n2988, Q => n10797, QN => n2519);
   REGISTERS_reg_76_23_inst : DFFR_X1 port map( D => n8757_port, CK => CLK, RN 
                           => n2987, Q => n10798, QN => n2520);
   REGISTERS_reg_76_22_inst : DFFR_X1 port map( D => n8758_port, CK => CLK, RN 
                           => n2987, Q => n10799, QN => n2521);
   REGISTERS_reg_76_21_inst : DFFR_X1 port map( D => n8759_port, CK => CLK, RN 
                           => n2987, Q => n10800, QN => n2522);
   REGISTERS_reg_76_20_inst : DFFR_X1 port map( D => n8760_port, CK => CLK, RN 
                           => n2987, Q => n10801, QN => n2523);
   REGISTERS_reg_76_19_inst : DFFR_X1 port map( D => n8761_port, CK => CLK, RN 
                           => n2987, Q => n10802, QN => n2524);
   REGISTERS_reg_76_18_inst : DFFR_X1 port map( D => n8762_port, CK => CLK, RN 
                           => n2987, Q => n10803, QN => n2525);
   REGISTERS_reg_76_17_inst : DFFR_X1 port map( D => n8763_port, CK => CLK, RN 
                           => n2987, Q => n10804, QN => n2526);
   REGISTERS_reg_76_16_inst : DFFR_X1 port map( D => n8764_port, CK => CLK, RN 
                           => n2987, Q => n10805, QN => n2527);
   REGISTERS_reg_76_15_inst : DFFR_X1 port map( D => n8765_port, CK => CLK, RN 
                           => n2987, Q => n10806, QN => n2528);
   REGISTERS_reg_76_14_inst : DFFR_X1 port map( D => n8766_port, CK => CLK, RN 
                           => n2987, Q => n10807, QN => n2529);
   REGISTERS_reg_76_13_inst : DFFR_X1 port map( D => n8767_port, CK => CLK, RN 
                           => n2987, Q => n10808, QN => n2530);
   REGISTERS_reg_76_12_inst : DFFR_X1 port map( D => n8768, CK => CLK, RN => 
                           n2987, Q => n10809, QN => n2531);
   REGISTERS_reg_76_11_inst : DFFR_X1 port map( D => n8769, CK => CLK, RN => 
                           n2986, Q => n10810, QN => n2532);
   REGISTERS_reg_76_10_inst : DFFR_X1 port map( D => n8770, CK => CLK, RN => 
                           n2986, Q => n10811, QN => n2533);
   REGISTERS_reg_76_9_inst : DFFR_X1 port map( D => n8771, CK => CLK, RN => 
                           n2986, Q => n10812, QN => n2534);
   REGISTERS_reg_76_8_inst : DFFR_X1 port map( D => n8772, CK => CLK, RN => 
                           n2986, Q => n10813, QN => n2535);
   REGISTERS_reg_76_7_inst : DFFR_X1 port map( D => n8773, CK => CLK, RN => 
                           n2986, Q => n10814, QN => n2536);
   REGISTERS_reg_76_6_inst : DFFR_X1 port map( D => n8774, CK => CLK, RN => 
                           n2986, Q => n10815, QN => n2537);
   REGISTERS_reg_76_5_inst : DFFR_X1 port map( D => n8775, CK => CLK, RN => 
                           n2986, Q => n10816, QN => n2538);
   REGISTERS_reg_76_4_inst : DFFR_X1 port map( D => n8776, CK => CLK, RN => 
                           n2986, Q => n10817, QN => n2539);
   REGISTERS_reg_76_3_inst : DFFR_X1 port map( D => n8777, CK => CLK, RN => 
                           n2986, Q => n10818, QN => n2540);
   REGISTERS_reg_76_2_inst : DFFR_X1 port map( D => n8778, CK => CLK, RN => 
                           n2986, Q => n10819, QN => n2541);
   REGISTERS_reg_76_1_inst : DFFR_X1 port map( D => n8779, CK => CLK, RN => 
                           n2986, Q => n10820, QN => n2542);
   REGISTERS_reg_76_0_inst : DFFR_X1 port map( D => n8780, CK => CLK, RN => 
                           n2986, Q => n10821, QN => n2543);
   REGISTERS_reg_79_31_inst : DFFR_X1 port map( D => n8845, CK => CLK, RN => 
                           n2980, Q => n10822, QN => n2608);
   REGISTERS_reg_79_30_inst : DFFR_X1 port map( D => n8846, CK => CLK, RN => 
                           n2980, Q => n10823, QN => n2609);
   REGISTERS_reg_79_29_inst : DFFR_X1 port map( D => n8847, CK => CLK, RN => 
                           n2980, Q => n10824, QN => n2610);
   REGISTERS_reg_79_28_inst : DFFR_X1 port map( D => n8848, CK => CLK, RN => 
                           n2980, Q => n10825, QN => n2611);
   REGISTERS_reg_79_27_inst : DFFR_X1 port map( D => n8849, CK => CLK, RN => 
                           n2980, Q => n10826, QN => n2612);
   REGISTERS_reg_79_26_inst : DFFR_X1 port map( D => n8850, CK => CLK, RN => 
                           n2980, Q => n10827, QN => n2613);
   REGISTERS_reg_79_25_inst : DFFR_X1 port map( D => n8851, CK => CLK, RN => 
                           n2980, Q => n10828, QN => n2614);
   REGISTERS_reg_79_24_inst : DFFR_X1 port map( D => n8852, CK => CLK, RN => 
                           n2980, Q => n10829, QN => n2615);
   REGISTERS_reg_79_23_inst : DFFR_X1 port map( D => n8853, CK => CLK, RN => 
                           n2979, Q => n10830, QN => n2616);
   REGISTERS_reg_79_22_inst : DFFR_X1 port map( D => n8854, CK => CLK, RN => 
                           n2979, Q => n10831, QN => n2617);
   REGISTERS_reg_79_21_inst : DFFR_X1 port map( D => n8855, CK => CLK, RN => 
                           n2979, Q => n10832, QN => n2618);
   REGISTERS_reg_79_20_inst : DFFR_X1 port map( D => n8856, CK => CLK, RN => 
                           n2979, Q => n10833, QN => n2619);
   REGISTERS_reg_79_19_inst : DFFR_X1 port map( D => n8857, CK => CLK, RN => 
                           n2979, Q => n10834, QN => n2620);
   REGISTERS_reg_79_18_inst : DFFR_X1 port map( D => n8858, CK => CLK, RN => 
                           n2979, Q => n10835, QN => n2621);
   REGISTERS_reg_79_17_inst : DFFR_X1 port map( D => n8859, CK => CLK, RN => 
                           n2979, Q => n10836, QN => n2622);
   REGISTERS_reg_79_16_inst : DFFR_X1 port map( D => n8860, CK => CLK, RN => 
                           n2979, Q => n10837, QN => n2623);
   REGISTERS_reg_79_15_inst : DFFR_X1 port map( D => n8861, CK => CLK, RN => 
                           n2979, Q => n10838, QN => n2624);
   REGISTERS_reg_79_14_inst : DFFR_X1 port map( D => n8862, CK => CLK, RN => 
                           n2979, Q => n10839, QN => n2625);
   REGISTERS_reg_79_13_inst : DFFR_X1 port map( D => n8863, CK => CLK, RN => 
                           n2979, Q => n10840, QN => n2626);
   REGISTERS_reg_79_12_inst : DFFR_X1 port map( D => n8864, CK => CLK, RN => 
                           n2979, Q => n10841, QN => n2627);
   REGISTERS_reg_79_11_inst : DFFR_X1 port map( D => n8865, CK => CLK, RN => 
                           n2978, Q => n10842, QN => n2628);
   REGISTERS_reg_79_10_inst : DFFR_X1 port map( D => n8866, CK => CLK, RN => 
                           n2978, Q => n10843, QN => n2629);
   REGISTERS_reg_79_9_inst : DFFR_X1 port map( D => n8867, CK => CLK, RN => 
                           n2978, Q => n10844, QN => n2630);
   REGISTERS_reg_79_8_inst : DFFR_X1 port map( D => n8868, CK => CLK, RN => 
                           n2978, Q => n10845, QN => n2631);
   REGISTERS_reg_79_7_inst : DFFR_X1 port map( D => n8869, CK => CLK, RN => 
                           n2978, Q => n10846, QN => n2632);
   REGISTERS_reg_79_6_inst : DFFR_X1 port map( D => n8870, CK => CLK, RN => 
                           n2978, Q => n10847, QN => n2633);
   REGISTERS_reg_79_5_inst : DFFR_X1 port map( D => n8871, CK => CLK, RN => 
                           n2978, Q => n10848, QN => n2634);
   REGISTERS_reg_79_4_inst : DFFR_X1 port map( D => n8872, CK => CLK, RN => 
                           n2978, Q => n10849, QN => n2635);
   REGISTERS_reg_79_3_inst : DFFR_X1 port map( D => n8873, CK => CLK, RN => 
                           n2978, Q => n10850, QN => n2636);
   REGISTERS_reg_79_2_inst : DFFR_X1 port map( D => n8874, CK => CLK, RN => 
                           n2978, Q => n10851, QN => n2637);
   REGISTERS_reg_79_1_inst : DFFR_X1 port map( D => n8875, CK => CLK, RN => 
                           n2978, Q => n10852, QN => n2638);
   REGISTERS_reg_79_0_inst : DFFR_X1 port map( D => n8876, CK => CLK, RN => 
                           n2978, Q => n10853, QN => n2639);
   REGISTERS_reg_80_31_inst : DFFR_X1 port map( D => n8877, CK => CLK, RN => 
                           n2977, Q => n10854, QN => n2640);
   REGISTERS_reg_80_30_inst : DFFR_X1 port map( D => n8878, CK => CLK, RN => 
                           n2977, Q => n10855, QN => n2641);
   REGISTERS_reg_80_29_inst : DFFR_X1 port map( D => n8879, CK => CLK, RN => 
                           n2977, Q => n10856, QN => n2642);
   REGISTERS_reg_80_28_inst : DFFR_X1 port map( D => n8880, CK => CLK, RN => 
                           n2977, Q => n10857, QN => n2643);
   REGISTERS_reg_80_27_inst : DFFR_X1 port map( D => n8881, CK => CLK, RN => 
                           n2977, Q => n10858, QN => n2644);
   REGISTERS_reg_80_26_inst : DFFR_X1 port map( D => n8882, CK => CLK, RN => 
                           n2977, Q => n10859, QN => n2645);
   REGISTERS_reg_80_25_inst : DFFR_X1 port map( D => n8883, CK => CLK, RN => 
                           n2977, Q => n10860, QN => n2646);
   REGISTERS_reg_80_24_inst : DFFR_X1 port map( D => n8884, CK => CLK, RN => 
                           n2977, Q => n10861, QN => n2647);
   REGISTERS_reg_80_23_inst : DFFR_X1 port map( D => n8885, CK => CLK, RN => 
                           n2977, Q => n10862, QN => n2648);
   REGISTERS_reg_80_22_inst : DFFR_X1 port map( D => n8886, CK => CLK, RN => 
                           n2977, Q => n10863, QN => n2649);
   REGISTERS_reg_80_21_inst : DFFR_X1 port map( D => n8887, CK => CLK, RN => 
                           n2977, Q => n10864, QN => n2650);
   REGISTERS_reg_80_20_inst : DFFR_X1 port map( D => n8888, CK => CLK, RN => 
                           n2977, Q => n10865, QN => n2651);
   REGISTERS_reg_80_19_inst : DFFR_X1 port map( D => n8889, CK => CLK, RN => 
                           n2976, Q => n10866, QN => n2652);
   REGISTERS_reg_80_18_inst : DFFR_X1 port map( D => n8890, CK => CLK, RN => 
                           n2976, Q => n10867, QN => n2653);
   REGISTERS_reg_80_17_inst : DFFR_X1 port map( D => n8891, CK => CLK, RN => 
                           n2976, Q => n10868, QN => n2654);
   REGISTERS_reg_80_16_inst : DFFR_X1 port map( D => n8892, CK => CLK, RN => 
                           n2976, Q => n10869, QN => n2655);
   REGISTERS_reg_80_15_inst : DFFR_X1 port map( D => n8893, CK => CLK, RN => 
                           n2976, Q => n10870, QN => n2656);
   REGISTERS_reg_80_14_inst : DFFR_X1 port map( D => n8894, CK => CLK, RN => 
                           n2976, Q => n10871, QN => n2657);
   REGISTERS_reg_80_13_inst : DFFR_X1 port map( D => n8895, CK => CLK, RN => 
                           n2976, Q => n10872, QN => n2658);
   REGISTERS_reg_80_12_inst : DFFR_X1 port map( D => n8896, CK => CLK, RN => 
                           n2976, Q => n10873, QN => n2659);
   REGISTERS_reg_80_11_inst : DFFR_X1 port map( D => n8897, CK => CLK, RN => 
                           n2976, Q => n10874, QN => n2660);
   REGISTERS_reg_80_10_inst : DFFR_X1 port map( D => n8898, CK => CLK, RN => 
                           n2976, Q => n10875, QN => n2661);
   REGISTERS_reg_80_9_inst : DFFR_X1 port map( D => n8899, CK => CLK, RN => 
                           n2976, Q => n10876, QN => n2662);
   REGISTERS_reg_80_8_inst : DFFR_X1 port map( D => n8900, CK => CLK, RN => 
                           n2976, Q => n10877, QN => n2663);
   REGISTERS_reg_80_7_inst : DFFR_X1 port map( D => n8901, CK => CLK, RN => 
                           n2975, Q => n10878, QN => n2664);
   REGISTERS_reg_80_6_inst : DFFR_X1 port map( D => n8902, CK => CLK, RN => 
                           n2975, Q => n10879, QN => n2665);
   REGISTERS_reg_80_5_inst : DFFR_X1 port map( D => n8903, CK => CLK, RN => 
                           n2975, Q => n10880, QN => n2666);
   REGISTERS_reg_80_4_inst : DFFR_X1 port map( D => n8904, CK => CLK, RN => 
                           n2975, Q => n10881, QN => n2667);
   REGISTERS_reg_80_3_inst : DFFR_X1 port map( D => n8905, CK => CLK, RN => 
                           n2975, Q => n10882, QN => n2668);
   REGISTERS_reg_80_2_inst : DFFR_X1 port map( D => n8906, CK => CLK, RN => 
                           n2975, Q => n10883, QN => n2669);
   REGISTERS_reg_80_1_inst : DFFR_X1 port map( D => n8907, CK => CLK, RN => 
                           n2975, Q => n10884, QN => n2670);
   REGISTERS_reg_80_0_inst : DFFR_X1 port map( D => n8908, CK => CLK, RN => 
                           n2975, Q => n10885, QN => n2671);
   REGISTERS_reg_81_31_inst : DFFR_X1 port map( D => n8909, CK => CLK, RN => 
                           n2975, Q => n10886, QN => n2672);
   REGISTERS_reg_81_30_inst : DFFR_X1 port map( D => n8910, CK => CLK, RN => 
                           n2975, Q => n10887, QN => n2673);
   REGISTERS_reg_81_29_inst : DFFR_X1 port map( D => n8911, CK => CLK, RN => 
                           n2975, Q => n10888, QN => n2674);
   REGISTERS_reg_81_28_inst : DFFR_X1 port map( D => n8912, CK => CLK, RN => 
                           n2975, Q => n10889, QN => n2675);
   REGISTERS_reg_81_27_inst : DFFR_X1 port map( D => n8913, CK => CLK, RN => 
                           n2974, Q => n10890, QN => n2676);
   REGISTERS_reg_81_26_inst : DFFR_X1 port map( D => n8914, CK => CLK, RN => 
                           n2974, Q => n10891, QN => n2677);
   REGISTERS_reg_81_25_inst : DFFR_X1 port map( D => n8915, CK => CLK, RN => 
                           n2974, Q => n10892, QN => n2678);
   REGISTERS_reg_81_24_inst : DFFR_X1 port map( D => n8916, CK => CLK, RN => 
                           n2974, Q => n10893, QN => n2679);
   REGISTERS_reg_81_23_inst : DFFR_X1 port map( D => n8917, CK => CLK, RN => 
                           n2974, Q => n10894, QN => n2680);
   REGISTERS_reg_81_22_inst : DFFR_X1 port map( D => n8918, CK => CLK, RN => 
                           n2974, Q => n10895, QN => n2681);
   REGISTERS_reg_81_21_inst : DFFR_X1 port map( D => n8919, CK => CLK, RN => 
                           n2974, Q => n10896, QN => n2682);
   REGISTERS_reg_81_20_inst : DFFR_X1 port map( D => n8920, CK => CLK, RN => 
                           n2974, Q => n10897, QN => n2683);
   REGISTERS_reg_81_19_inst : DFFR_X1 port map( D => n8921, CK => CLK, RN => 
                           n2974, Q => n10898, QN => n2684);
   REGISTERS_reg_81_18_inst : DFFR_X1 port map( D => n8922, CK => CLK, RN => 
                           n2974, Q => n10899, QN => n2685);
   REGISTERS_reg_81_17_inst : DFFR_X1 port map( D => n8923, CK => CLK, RN => 
                           n2974, Q => n10900, QN => n2686);
   REGISTERS_reg_81_16_inst : DFFR_X1 port map( D => n8924, CK => CLK, RN => 
                           n2974, Q => n10901, QN => n2687);
   REGISTERS_reg_81_15_inst : DFFR_X1 port map( D => n8925, CK => CLK, RN => 
                           n2973, Q => n10902, QN => n2688);
   REGISTERS_reg_81_14_inst : DFFR_X1 port map( D => n8926, CK => CLK, RN => 
                           n2973, Q => n10903, QN => n2689);
   REGISTERS_reg_81_13_inst : DFFR_X1 port map( D => n8927, CK => CLK, RN => 
                           n2973, Q => n10904, QN => n2690);
   REGISTERS_reg_81_12_inst : DFFR_X1 port map( D => n8928, CK => CLK, RN => 
                           n2973, Q => n10905, QN => n2691);
   REGISTERS_reg_81_11_inst : DFFR_X1 port map( D => n8929, CK => CLK, RN => 
                           n2973, Q => n10906, QN => n2692);
   REGISTERS_reg_81_10_inst : DFFR_X1 port map( D => n8930, CK => CLK, RN => 
                           n2973, Q => n10907, QN => n2693);
   REGISTERS_reg_81_9_inst : DFFR_X1 port map( D => n8931, CK => CLK, RN => 
                           n2973, Q => n10908, QN => n2694);
   REGISTERS_reg_81_8_inst : DFFR_X1 port map( D => n8932, CK => CLK, RN => 
                           n2973, Q => n10909, QN => n2695);
   REGISTERS_reg_81_7_inst : DFFR_X1 port map( D => n8933, CK => CLK, RN => 
                           n2973, Q => n10910, QN => n2696);
   REGISTERS_reg_81_6_inst : DFFR_X1 port map( D => n8934, CK => CLK, RN => 
                           n2973, Q => n10911, QN => n2697);
   REGISTERS_reg_81_5_inst : DFFR_X1 port map( D => n8935, CK => CLK, RN => 
                           n2973, Q => n10912, QN => n2698);
   REGISTERS_reg_81_4_inst : DFFR_X1 port map( D => n8936, CK => CLK, RN => 
                           n2973, Q => n10913, QN => n2699);
   REGISTERS_reg_81_3_inst : DFFR_X1 port map( D => n8937, CK => CLK, RN => 
                           n2972, Q => n10914, QN => n2700);
   REGISTERS_reg_81_2_inst : DFFR_X1 port map( D => n8938, CK => CLK, RN => 
                           n2972, Q => n10915, QN => n2701);
   REGISTERS_reg_81_1_inst : DFFR_X1 port map( D => n8939, CK => CLK, RN => 
                           n2972, Q => n10916, QN => n2702);
   REGISTERS_reg_81_0_inst : DFFR_X1 port map( D => n8940, CK => CLK, RN => 
                           n2972, Q => n10917, QN => n2703);
   OUT2_reg_31_inst : DLH_X1 port map( G => n1791, D => N8767, Q => OUT2(31));
   OUT1_reg_31_inst : DLH_X1 port map( G => n1794, D => N8734, Q => OUT1(31));
   OUT2_reg_30_inst : DLH_X1 port map( G => n1791, D => N8766, Q => OUT2(30));
   OUT1_reg_30_inst : DLH_X1 port map( G => n1794, D => N8733, Q => OUT1(30));
   OUT2_reg_29_inst : DLH_X1 port map( G => n1791, D => N8765, Q => OUT2(29));
   OUT1_reg_29_inst : DLH_X1 port map( G => n1794, D => N8732, Q => OUT1(29));
   OUT2_reg_28_inst : DLH_X1 port map( G => n1791, D => N8764, Q => OUT2(28));
   OUT1_reg_28_inst : DLH_X1 port map( G => n1794, D => N8731, Q => OUT1(28));
   OUT2_reg_27_inst : DLH_X1 port map( G => n1791, D => N8763, Q => OUT2(27));
   OUT1_reg_27_inst : DLH_X1 port map( G => n1794, D => N8730, Q => OUT1(27));
   OUT2_reg_26_inst : DLH_X1 port map( G => n1791, D => N8762, Q => OUT2(26));
   OUT1_reg_26_inst : DLH_X1 port map( G => n1794, D => N8729, Q => OUT1(26));
   OUT2_reg_25_inst : DLH_X1 port map( G => n1791, D => N8761, Q => OUT2(25));
   OUT1_reg_25_inst : DLH_X1 port map( G => n1794, D => N8728, Q => OUT1(25));
   OUT2_reg_24_inst : DLH_X1 port map( G => n1791, D => N8760, Q => OUT2(24));
   OUT1_reg_24_inst : DLH_X1 port map( G => n1794, D => N8727, Q => OUT1(24));
   OUT2_reg_23_inst : DLH_X1 port map( G => n1791, D => N8759, Q => OUT2(23));
   OUT1_reg_23_inst : DLH_X1 port map( G => n1794, D => N8726, Q => OUT1(23));
   OUT2_reg_22_inst : DLH_X1 port map( G => n1791, D => N8758, Q => OUT2(22));
   OUT1_reg_22_inst : DLH_X1 port map( G => n1794, D => N8725, Q => OUT1(22));
   OUT2_reg_21_inst : DLH_X1 port map( G => n1791, D => N8757, Q => OUT2(21));
   OUT1_reg_21_inst : DLH_X1 port map( G => n1794, D => N8724, Q => OUT1(21));
   OUT2_reg_20_inst : DLH_X1 port map( G => n1792, D => N8756, Q => OUT2(20));
   OUT1_reg_20_inst : DLH_X1 port map( G => n1795, D => N8723, Q => OUT1(20));
   OUT2_reg_19_inst : DLH_X1 port map( G => n1792, D => N8755, Q => OUT2(19));
   OUT1_reg_19_inst : DLH_X1 port map( G => n1795, D => N8722, Q => OUT1(19));
   OUT2_reg_18_inst : DLH_X1 port map( G => n1792, D => N8754, Q => OUT2(18));
   OUT1_reg_18_inst : DLH_X1 port map( G => n1795, D => N8721, Q => OUT1(18));
   OUT2_reg_17_inst : DLH_X1 port map( G => n1792, D => N8753, Q => OUT2(17));
   OUT1_reg_17_inst : DLH_X1 port map( G => n1795, D => N8720, Q => OUT1(17));
   OUT2_reg_16_inst : DLH_X1 port map( G => n1792, D => N8752, Q => OUT2(16));
   OUT1_reg_16_inst : DLH_X1 port map( G => n1795, D => N8719, Q => OUT1(16));
   OUT2_reg_15_inst : DLH_X1 port map( G => n1792, D => N8751, Q => OUT2(15));
   OUT1_reg_15_inst : DLH_X1 port map( G => n1795, D => N8718, Q => OUT1(15));
   OUT2_reg_14_inst : DLH_X1 port map( G => n1792, D => N8750, Q => OUT2(14));
   OUT1_reg_14_inst : DLH_X1 port map( G => n1795, D => N8717, Q => OUT1(14));
   OUT2_reg_13_inst : DLH_X1 port map( G => n1792, D => N8749, Q => OUT2(13));
   OUT1_reg_13_inst : DLH_X1 port map( G => n1795, D => N8716, Q => OUT1(13));
   OUT2_reg_12_inst : DLH_X1 port map( G => n1792, D => N8748, Q => OUT2(12));
   OUT1_reg_12_inst : DLH_X1 port map( G => n1795, D => N8715, Q => OUT1(12));
   OUT2_reg_11_inst : DLH_X1 port map( G => n1792, D => N8747, Q => OUT2(11));
   OUT1_reg_11_inst : DLH_X1 port map( G => n1795, D => N8714, Q => OUT1(11));
   OUT2_reg_10_inst : DLH_X1 port map( G => n1792, D => N8746, Q => OUT2(10));
   OUT1_reg_10_inst : DLH_X1 port map( G => n1795, D => N8713, Q => OUT1(10));
   OUT2_reg_9_inst : DLH_X1 port map( G => n1793, D => N8745, Q => OUT2(9));
   OUT1_reg_9_inst : DLH_X1 port map( G => n1796, D => N8712, Q => OUT1(9));
   OUT2_reg_8_inst : DLH_X1 port map( G => n1793, D => N8744, Q => OUT2(8));
   OUT1_reg_8_inst : DLH_X1 port map( G => n1796, D => N8711, Q => OUT1(8));
   OUT2_reg_7_inst : DLH_X1 port map( G => n1793, D => N8743, Q => OUT2(7));
   OUT1_reg_7_inst : DLH_X1 port map( G => n1796, D => N8710, Q => OUT1(7));
   OUT2_reg_6_inst : DLH_X1 port map( G => n1793, D => N8742, Q => OUT2(6));
   OUT1_reg_6_inst : DLH_X1 port map( G => n1796, D => N8709, Q => OUT1(6));
   OUT2_reg_5_inst : DLH_X1 port map( G => n1793, D => N8741, Q => OUT2(5));
   OUT1_reg_5_inst : DLH_X1 port map( G => n1796, D => N8708, Q => OUT1(5));
   OUT2_reg_4_inst : DLH_X1 port map( G => n1793, D => N8740, Q => OUT2(4));
   OUT1_reg_4_inst : DLH_X1 port map( G => n1796, D => N8707, Q => OUT1(4));
   OUT2_reg_3_inst : DLH_X1 port map( G => n1793, D => N8739, Q => OUT2(3));
   OUT1_reg_3_inst : DLH_X1 port map( G => n1796, D => N8706, Q => OUT1(3));
   OUT2_reg_2_inst : DLH_X1 port map( G => n1793, D => N8738, Q => OUT2(2));
   OUT1_reg_2_inst : DLH_X1 port map( G => n1796, D => N8705, Q => OUT1(2));
   OUT2_reg_1_inst : DLH_X1 port map( G => n1793, D => N8737, Q => OUT2(1));
   OUT1_reg_1_inst : DLH_X1 port map( G => n1796, D => N8704, Q => OUT1(1));
   OUT2_reg_0_inst : DLH_X1 port map( G => n1793, D => N8736, Q => OUT2(0));
   OUT1_reg_0_inst : DLH_X1 port map( G => n1796, D => N8703, Q => OUT1(0));
   FILL <= '0';
   SPILL <= '0';
   add_66_C130 : windRF_M8_N8_F5_NBIT32_DW01_add_1 port map( A(6) => CWP_6_port
                           , A(5) => CWP_5_port, A(4) => CWP_4_port, A(3) => 
                           N8790, A(2) => N8789, A(1) => N8788, A(0) => N8787, 
                           B(6) => n7, B(5) => n7, B(4) => ADD_RD2(4), B(3) => 
                           ADD_RD2(3), B(2) => ADD_RD2(2), B(1) => ADD_RD2(1), 
                           B(0) => ADD_RD2(0), CI => n7, SUM(6) => N8567, 
                           SUM(5) => N8566, SUM(4) => N8565, SUM(3) => N8564, 
                           SUM(2) => N8563, SUM(1) => N8562, SUM(0) => N8561, 
                           CO => n_1185);
   add_66_C126 : windRF_M8_N8_F5_NBIT32_DW01_add_3 port map( A(6) => CWP_6_port
                           , A(5) => CWP_5_port, A(4) => CWP_4_port, A(3) => 
                           N8790, A(2) => N8789, A(1) => N8788, A(0) => N8787, 
                           B(6) => n11, B(5) => n11, B(4) => ADD_RD1(4), B(3) 
                           => ADD_RD1(3), B(2) => ADD_RD1(2), B(1) => 
                           ADD_RD1(1), B(0) => ADD_RD1(0), CI => n11, SUM(6) =>
                           N8423, SUM(5) => N8422, SUM(4) => N8421, SUM(3) => 
                           N8420, SUM(2) => N8419, SUM(1) => N8418, SUM(0) => 
                           N8417, CO => n_1186);
   add_66_C91 : windRF_M8_N8_F5_NBIT32_DW01_add_5 port map( A(6) => CWP_6_port,
                           A(5) => CWP_5_port, A(4) => CWP_4_port, A(3) => 
                           N8790, A(2) => N8789, A(1) => N8788, A(0) => N8787, 
                           B(6) => n17, B(5) => n17, B(4) => ADD_WR(4), B(3) =>
                           ADD_WR(3), B(2) => ADD_WR(2), B(1) => ADD_WR(1), 
                           B(0) => ADD_WR(0), CI => n17, SUM(6) => N2159, 
                           SUM(5) => N2158, SUM(4) => N2157, SUM(3) => N2156, 
                           SUM(2) => N2155, SUM(1) => N2154, SUM(0) => N2153, 
                           CO => n_1187);
   REGISTERS_reg_87_31_inst : DFFR_X1 port map( D => n9101, CK => CLK, RN => 
                           RESET, Q => REGISTERS_87_31_port, QN => n_1188);
   REGISTERS_reg_87_30_inst : DFFR_X1 port map( D => n9102, CK => CLK, RN => 
                           n2959, Q => REGISTERS_87_30_port, QN => n_1189);
   REGISTERS_reg_87_29_inst : DFFR_X1 port map( D => n9103, CK => CLK, RN => 
                           n2959, Q => REGISTERS_87_29_port, QN => n_1190);
   REGISTERS_reg_87_28_inst : DFFR_X1 port map( D => n9104, CK => CLK, RN => 
                           n2959, Q => REGISTERS_87_28_port, QN => n_1191);
   REGISTERS_reg_87_27_inst : DFFR_X1 port map( D => n9105, CK => CLK, RN => 
                           n2958, Q => REGISTERS_87_27_port, QN => n_1192);
   REGISTERS_reg_87_26_inst : DFFR_X1 port map( D => n9106, CK => CLK, RN => 
                           n2958, Q => REGISTERS_87_26_port, QN => n_1193);
   REGISTERS_reg_87_25_inst : DFFR_X1 port map( D => n9107, CK => CLK, RN => 
                           n2958, Q => REGISTERS_87_25_port, QN => n_1194);
   REGISTERS_reg_87_24_inst : DFFR_X1 port map( D => n9108, CK => CLK, RN => 
                           n2958, Q => REGISTERS_87_24_port, QN => n_1195);
   REGISTERS_reg_87_23_inst : DFFR_X1 port map( D => n9109, CK => CLK, RN => 
                           n2958, Q => REGISTERS_87_23_port, QN => n_1196);
   REGISTERS_reg_87_22_inst : DFFR_X1 port map( D => n9110, CK => CLK, RN => 
                           n2958, Q => REGISTERS_87_22_port, QN => n_1197);
   REGISTERS_reg_87_21_inst : DFFR_X1 port map( D => n9111, CK => CLK, RN => 
                           n2958, Q => REGISTERS_87_21_port, QN => n_1198);
   REGISTERS_reg_87_20_inst : DFFR_X1 port map( D => n9112, CK => CLK, RN => 
                           n2958, Q => REGISTERS_87_20_port, QN => n_1199);
   REGISTERS_reg_87_19_inst : DFFR_X1 port map( D => n9113, CK => CLK, RN => 
                           n2958, Q => REGISTERS_87_19_port, QN => n_1200);
   REGISTERS_reg_87_18_inst : DFFR_X1 port map( D => n9114, CK => CLK, RN => 
                           n2958, Q => REGISTERS_87_18_port, QN => n_1201);
   REGISTERS_reg_87_17_inst : DFFR_X1 port map( D => n9115, CK => CLK, RN => 
                           n2958, Q => REGISTERS_87_17_port, QN => n_1202);
   REGISTERS_reg_87_16_inst : DFFR_X1 port map( D => n9116, CK => CLK, RN => 
                           n2958, Q => REGISTERS_87_16_port, QN => n_1203);
   REGISTERS_reg_87_15_inst : DFFR_X1 port map( D => n9117, CK => CLK, RN => 
                           n2957, Q => REGISTERS_87_15_port, QN => n_1204);
   REGISTERS_reg_87_14_inst : DFFR_X1 port map( D => n9118, CK => CLK, RN => 
                           n2957, Q => REGISTERS_87_14_port, QN => n_1205);
   REGISTERS_reg_87_13_inst : DFFR_X1 port map( D => n9119, CK => CLK, RN => 
                           n2957, Q => REGISTERS_87_13_port, QN => n_1206);
   REGISTERS_reg_87_12_inst : DFFR_X1 port map( D => n9120, CK => CLK, RN => 
                           n2957, Q => REGISTERS_87_12_port, QN => n_1207);
   REGISTERS_reg_87_11_inst : DFFR_X1 port map( D => n9121, CK => CLK, RN => 
                           n2957, Q => REGISTERS_87_11_port, QN => n_1208);
   REGISTERS_reg_87_10_inst : DFFR_X1 port map( D => n9122, CK => CLK, RN => 
                           n2957, Q => REGISTERS_87_10_port, QN => n_1209);
   REGISTERS_reg_87_9_inst : DFFR_X1 port map( D => n9123, CK => CLK, RN => 
                           n2957, Q => REGISTERS_87_9_port, QN => n_1210);
   REGISTERS_reg_87_8_inst : DFFR_X1 port map( D => n9124, CK => CLK, RN => 
                           n2957, Q => REGISTERS_87_8_port, QN => n_1211);
   REGISTERS_reg_87_7_inst : DFFR_X1 port map( D => n9125, CK => CLK, RN => 
                           n2957, Q => REGISTERS_87_7_port, QN => n_1212);
   REGISTERS_reg_87_6_inst : DFFR_X1 port map( D => n9126, CK => CLK, RN => 
                           n2957, Q => REGISTERS_87_6_port, QN => n_1213);
   REGISTERS_reg_87_5_inst : DFFR_X1 port map( D => n9127, CK => CLK, RN => 
                           n2957, Q => REGISTERS_87_5_port, QN => n_1214);
   REGISTERS_reg_87_4_inst : DFFR_X1 port map( D => n9128, CK => CLK, RN => 
                           n2957, Q => REGISTERS_87_4_port, QN => n_1215);
   REGISTERS_reg_87_3_inst : DFFR_X1 port map( D => n9129, CK => CLK, RN => 
                           n2956, Q => REGISTERS_87_3_port, QN => n_1216);
   REGISTERS_reg_87_2_inst : DFFR_X1 port map( D => n9130, CK => CLK, RN => 
                           n2956, Q => REGISTERS_87_2_port, QN => n_1217);
   REGISTERS_reg_87_1_inst : DFFR_X1 port map( D => n9131, CK => CLK, RN => 
                           n2956, Q => REGISTERS_87_1_port, QN => n_1218);
   REGISTERS_reg_87_0_inst : DFFR_X1 port map( D => n9132, CK => CLK, RN => 
                           n2956, Q => REGISTERS_87_0_port, QN => n_1219);
   REGISTERS_reg_86_31_inst : DFFR_X1 port map( D => n9069, CK => CLK, RN => 
                           n2961, Q => REGISTERS_86_31_port, QN => n_1220);
   REGISTERS_reg_86_30_inst : DFFR_X1 port map( D => n9070, CK => CLK, RN => 
                           n2961, Q => REGISTERS_86_30_port, QN => n_1221);
   REGISTERS_reg_86_29_inst : DFFR_X1 port map( D => n9071, CK => CLK, RN => 
                           n2961, Q => REGISTERS_86_29_port, QN => n_1222);
   REGISTERS_reg_86_28_inst : DFFR_X1 port map( D => n9072, CK => CLK, RN => 
                           n2961, Q => REGISTERS_86_28_port, QN => n_1223);
   REGISTERS_reg_86_27_inst : DFFR_X1 port map( D => n9073, CK => CLK, RN => 
                           n2961, Q => REGISTERS_86_27_port, QN => n_1224);
   REGISTERS_reg_86_26_inst : DFFR_X1 port map( D => n9074, CK => CLK, RN => 
                           n2961, Q => REGISTERS_86_26_port, QN => n_1225);
   REGISTERS_reg_86_25_inst : DFFR_X1 port map( D => n9075, CK => CLK, RN => 
                           n2961, Q => REGISTERS_86_25_port, QN => n_1226);
   REGISTERS_reg_86_24_inst : DFFR_X1 port map( D => n9076, CK => CLK, RN => 
                           n2961, Q => REGISTERS_86_24_port, QN => n_1227);
   REGISTERS_reg_86_23_inst : DFFR_X1 port map( D => n9077, CK => CLK, RN => 
                           n2961, Q => REGISTERS_86_23_port, QN => n_1228);
   REGISTERS_reg_86_22_inst : DFFR_X1 port map( D => n9078, CK => CLK, RN => 
                           n2961, Q => REGISTERS_86_22_port, QN => n_1229);
   REGISTERS_reg_86_21_inst : DFFR_X1 port map( D => n9079, CK => CLK, RN => 
                           n2961, Q => REGISTERS_86_21_port, QN => n_1230);
   REGISTERS_reg_86_20_inst : DFFR_X1 port map( D => n9080, CK => CLK, RN => 
                           n2961, Q => REGISTERS_86_20_port, QN => n_1231);
   REGISTERS_reg_86_19_inst : DFFR_X1 port map( D => n9081, CK => CLK, RN => 
                           n2960, Q => REGISTERS_86_19_port, QN => n_1232);
   REGISTERS_reg_86_18_inst : DFFR_X1 port map( D => n9082, CK => CLK, RN => 
                           n2960, Q => REGISTERS_86_18_port, QN => n_1233);
   REGISTERS_reg_86_17_inst : DFFR_X1 port map( D => n9083, CK => CLK, RN => 
                           n2960, Q => REGISTERS_86_17_port, QN => n_1234);
   REGISTERS_reg_86_16_inst : DFFR_X1 port map( D => n9084, CK => CLK, RN => 
                           n2960, Q => REGISTERS_86_16_port, QN => n_1235);
   REGISTERS_reg_86_15_inst : DFFR_X1 port map( D => n9085, CK => CLK, RN => 
                           n2960, Q => REGISTERS_86_15_port, QN => n_1236);
   REGISTERS_reg_86_14_inst : DFFR_X1 port map( D => n9086, CK => CLK, RN => 
                           n2960, Q => REGISTERS_86_14_port, QN => n_1237);
   REGISTERS_reg_86_13_inst : DFFR_X1 port map( D => n9087, CK => CLK, RN => 
                           n2960, Q => REGISTERS_86_13_port, QN => n_1238);
   REGISTERS_reg_86_12_inst : DFFR_X1 port map( D => n9088, CK => CLK, RN => 
                           n2960, Q => REGISTERS_86_12_port, QN => n_1239);
   REGISTERS_reg_86_11_inst : DFFR_X1 port map( D => n9089, CK => CLK, RN => 
                           n2960, Q => REGISTERS_86_11_port, QN => n_1240);
   REGISTERS_reg_86_10_inst : DFFR_X1 port map( D => n9090, CK => CLK, RN => 
                           n2960, Q => REGISTERS_86_10_port, QN => n_1241);
   REGISTERS_reg_86_9_inst : DFFR_X1 port map( D => n9091, CK => CLK, RN => 
                           n2960, Q => REGISTERS_86_9_port, QN => n_1242);
   REGISTERS_reg_86_8_inst : DFFR_X1 port map( D => n9092, CK => CLK, RN => 
                           n2960, Q => REGISTERS_86_8_port, QN => n_1243);
   REGISTERS_reg_86_7_inst : DFFR_X1 port map( D => n9093, CK => CLK, RN => 
                           n2959, Q => REGISTERS_86_7_port, QN => n_1244);
   REGISTERS_reg_86_6_inst : DFFR_X1 port map( D => n9094, CK => CLK, RN => 
                           n2959, Q => REGISTERS_86_6_port, QN => n_1245);
   REGISTERS_reg_86_5_inst : DFFR_X1 port map( D => n9095, CK => CLK, RN => 
                           n2959, Q => REGISTERS_86_5_port, QN => n_1246);
   REGISTERS_reg_86_4_inst : DFFR_X1 port map( D => n9096, CK => CLK, RN => 
                           n2959, Q => REGISTERS_86_4_port, QN => n_1247);
   REGISTERS_reg_86_3_inst : DFFR_X1 port map( D => n9097, CK => CLK, RN => 
                           n2959, Q => REGISTERS_86_3_port, QN => n_1248);
   REGISTERS_reg_86_2_inst : DFFR_X1 port map( D => n9098, CK => CLK, RN => 
                           n2959, Q => REGISTERS_86_2_port, QN => n_1249);
   REGISTERS_reg_86_1_inst : DFFR_X1 port map( D => n9099, CK => CLK, RN => 
                           n2959, Q => REGISTERS_86_1_port, QN => n_1250);
   REGISTERS_reg_86_0_inst : DFFR_X1 port map( D => n9100, CK => CLK, RN => 
                           n2959, Q => REGISTERS_86_0_port, QN => n_1251);
   REGISTERS_reg_85_31_inst : DFFR_X1 port map( D => n9037, CK => CLK, RN => 
                           n2964, Q => REGISTERS_85_31_port, QN => n_1252);
   REGISTERS_reg_85_30_inst : DFFR_X1 port map( D => n9038, CK => CLK, RN => 
                           n2964, Q => REGISTERS_85_30_port, QN => n_1253);
   REGISTERS_reg_85_29_inst : DFFR_X1 port map( D => n9039, CK => CLK, RN => 
                           n2964, Q => REGISTERS_85_29_port, QN => n_1254);
   REGISTERS_reg_85_28_inst : DFFR_X1 port map( D => n9040, CK => CLK, RN => 
                           n2964, Q => REGISTERS_85_28_port, QN => n_1255);
   REGISTERS_reg_85_27_inst : DFFR_X1 port map( D => n9041, CK => CLK, RN => 
                           n2964, Q => REGISTERS_85_27_port, QN => n_1256);
   REGISTERS_reg_85_26_inst : DFFR_X1 port map( D => n9042, CK => CLK, RN => 
                           n2964, Q => REGISTERS_85_26_port, QN => n_1257);
   REGISTERS_reg_85_25_inst : DFFR_X1 port map( D => n9043, CK => CLK, RN => 
                           n2964, Q => REGISTERS_85_25_port, QN => n_1258);
   REGISTERS_reg_85_24_inst : DFFR_X1 port map( D => n9044, CK => CLK, RN => 
                           n2964, Q => REGISTERS_85_24_port, QN => n_1259);
   REGISTERS_reg_85_23_inst : DFFR_X1 port map( D => n9045, CK => CLK, RN => 
                           n2963, Q => REGISTERS_85_23_port, QN => n_1260);
   REGISTERS_reg_85_22_inst : DFFR_X1 port map( D => n9046, CK => CLK, RN => 
                           n2963, Q => REGISTERS_85_22_port, QN => n_1261);
   REGISTERS_reg_85_21_inst : DFFR_X1 port map( D => n9047, CK => CLK, RN => 
                           n2963, Q => REGISTERS_85_21_port, QN => n_1262);
   REGISTERS_reg_85_20_inst : DFFR_X1 port map( D => n9048, CK => CLK, RN => 
                           n2963, Q => REGISTERS_85_20_port, QN => n_1263);
   REGISTERS_reg_85_19_inst : DFFR_X1 port map( D => n9049, CK => CLK, RN => 
                           n2963, Q => REGISTERS_85_19_port, QN => n_1264);
   REGISTERS_reg_85_18_inst : DFFR_X1 port map( D => n9050, CK => CLK, RN => 
                           n2963, Q => REGISTERS_85_18_port, QN => n_1265);
   REGISTERS_reg_85_17_inst : DFFR_X1 port map( D => n9051, CK => CLK, RN => 
                           n2963, Q => REGISTERS_85_17_port, QN => n_1266);
   REGISTERS_reg_85_16_inst : DFFR_X1 port map( D => n9052, CK => CLK, RN => 
                           n2963, Q => REGISTERS_85_16_port, QN => n_1267);
   REGISTERS_reg_85_15_inst : DFFR_X1 port map( D => n9053, CK => CLK, RN => 
                           n2963, Q => REGISTERS_85_15_port, QN => n_1268);
   REGISTERS_reg_85_14_inst : DFFR_X1 port map( D => n9054, CK => CLK, RN => 
                           n2963, Q => REGISTERS_85_14_port, QN => n_1269);
   REGISTERS_reg_85_13_inst : DFFR_X1 port map( D => n9055, CK => CLK, RN => 
                           n2963, Q => REGISTERS_85_13_port, QN => n_1270);
   REGISTERS_reg_85_12_inst : DFFR_X1 port map( D => n9056, CK => CLK, RN => 
                           n2963, Q => REGISTERS_85_12_port, QN => n_1271);
   REGISTERS_reg_85_11_inst : DFFR_X1 port map( D => n9057, CK => CLK, RN => 
                           n2962, Q => REGISTERS_85_11_port, QN => n_1272);
   REGISTERS_reg_85_10_inst : DFFR_X1 port map( D => n9058, CK => CLK, RN => 
                           n2962, Q => REGISTERS_85_10_port, QN => n_1273);
   REGISTERS_reg_85_9_inst : DFFR_X1 port map( D => n9059, CK => CLK, RN => 
                           n2962, Q => REGISTERS_85_9_port, QN => n_1274);
   REGISTERS_reg_85_8_inst : DFFR_X1 port map( D => n9060, CK => CLK, RN => 
                           n2962, Q => REGISTERS_85_8_port, QN => n_1275);
   REGISTERS_reg_85_7_inst : DFFR_X1 port map( D => n9061, CK => CLK, RN => 
                           n2962, Q => REGISTERS_85_7_port, QN => n_1276);
   REGISTERS_reg_85_6_inst : DFFR_X1 port map( D => n9062, CK => CLK, RN => 
                           n2962, Q => REGISTERS_85_6_port, QN => n_1277);
   REGISTERS_reg_85_5_inst : DFFR_X1 port map( D => n9063, CK => CLK, RN => 
                           n2962, Q => REGISTERS_85_5_port, QN => n_1278);
   REGISTERS_reg_85_4_inst : DFFR_X1 port map( D => n9064, CK => CLK, RN => 
                           n2962, Q => REGISTERS_85_4_port, QN => n_1279);
   REGISTERS_reg_85_3_inst : DFFR_X1 port map( D => n9065, CK => CLK, RN => 
                           n2962, Q => REGISTERS_85_3_port, QN => n_1280);
   REGISTERS_reg_85_2_inst : DFFR_X1 port map( D => n9066, CK => CLK, RN => 
                           n2962, Q => REGISTERS_85_2_port, QN => n_1281);
   REGISTERS_reg_85_1_inst : DFFR_X1 port map( D => n9067, CK => CLK, RN => 
                           n2962, Q => REGISTERS_85_1_port, QN => n_1282);
   REGISTERS_reg_85_0_inst : DFFR_X1 port map( D => n9068, CK => CLK, RN => 
                           n2962, Q => REGISTERS_85_0_port, QN => n_1283);
   REGISTERS_reg_84_31_inst : DFFR_X1 port map( D => n9005, CK => CLK, RN => 
                           n2967, Q => REGISTERS_84_31_port, QN => n_1284);
   REGISTERS_reg_84_30_inst : DFFR_X1 port map( D => n9006, CK => CLK, RN => 
                           n2967, Q => REGISTERS_84_30_port, QN => n_1285);
   REGISTERS_reg_84_29_inst : DFFR_X1 port map( D => n9007, CK => CLK, RN => 
                           n2967, Q => REGISTERS_84_29_port, QN => n_1286);
   REGISTERS_reg_84_28_inst : DFFR_X1 port map( D => n9008, CK => CLK, RN => 
                           n2967, Q => REGISTERS_84_28_port, QN => n_1287);
   REGISTERS_reg_84_27_inst : DFFR_X1 port map( D => n9009, CK => CLK, RN => 
                           n2966, Q => REGISTERS_84_27_port, QN => n_1288);
   REGISTERS_reg_84_26_inst : DFFR_X1 port map( D => n9010, CK => CLK, RN => 
                           n2966, Q => REGISTERS_84_26_port, QN => n_1289);
   REGISTERS_reg_84_25_inst : DFFR_X1 port map( D => n9011, CK => CLK, RN => 
                           n2966, Q => REGISTERS_84_25_port, QN => n_1290);
   REGISTERS_reg_84_24_inst : DFFR_X1 port map( D => n9012, CK => CLK, RN => 
                           n2966, Q => REGISTERS_84_24_port, QN => n_1291);
   REGISTERS_reg_84_23_inst : DFFR_X1 port map( D => n9013, CK => CLK, RN => 
                           n2966, Q => REGISTERS_84_23_port, QN => n_1292);
   REGISTERS_reg_84_22_inst : DFFR_X1 port map( D => n9014, CK => CLK, RN => 
                           n2966, Q => REGISTERS_84_22_port, QN => n_1293);
   REGISTERS_reg_84_21_inst : DFFR_X1 port map( D => n9015, CK => CLK, RN => 
                           n2966, Q => REGISTERS_84_21_port, QN => n_1294);
   REGISTERS_reg_84_20_inst : DFFR_X1 port map( D => n9016, CK => CLK, RN => 
                           n2966, Q => REGISTERS_84_20_port, QN => n_1295);
   REGISTERS_reg_84_19_inst : DFFR_X1 port map( D => n9017, CK => CLK, RN => 
                           n2966, Q => REGISTERS_84_19_port, QN => n_1296);
   REGISTERS_reg_84_18_inst : DFFR_X1 port map( D => n9018, CK => CLK, RN => 
                           n2966, Q => REGISTERS_84_18_port, QN => n_1297);
   REGISTERS_reg_84_17_inst : DFFR_X1 port map( D => n9019, CK => CLK, RN => 
                           n2966, Q => REGISTERS_84_17_port, QN => n_1298);
   REGISTERS_reg_84_16_inst : DFFR_X1 port map( D => n9020, CK => CLK, RN => 
                           n2966, Q => REGISTERS_84_16_port, QN => n_1299);
   REGISTERS_reg_84_15_inst : DFFR_X1 port map( D => n9021, CK => CLK, RN => 
                           n2965, Q => REGISTERS_84_15_port, QN => n_1300);
   REGISTERS_reg_84_14_inst : DFFR_X1 port map( D => n9022, CK => CLK, RN => 
                           n2965, Q => REGISTERS_84_14_port, QN => n_1301);
   REGISTERS_reg_84_13_inst : DFFR_X1 port map( D => n9023, CK => CLK, RN => 
                           n2965, Q => REGISTERS_84_13_port, QN => n_1302);
   REGISTERS_reg_84_12_inst : DFFR_X1 port map( D => n9024, CK => CLK, RN => 
                           n2965, Q => REGISTERS_84_12_port, QN => n_1303);
   REGISTERS_reg_84_11_inst : DFFR_X1 port map( D => n9025, CK => CLK, RN => 
                           n2965, Q => REGISTERS_84_11_port, QN => n_1304);
   REGISTERS_reg_84_10_inst : DFFR_X1 port map( D => n9026, CK => CLK, RN => 
                           n2965, Q => REGISTERS_84_10_port, QN => n_1305);
   REGISTERS_reg_84_9_inst : DFFR_X1 port map( D => n9027, CK => CLK, RN => 
                           n2965, Q => REGISTERS_84_9_port, QN => n_1306);
   REGISTERS_reg_84_8_inst : DFFR_X1 port map( D => n9028, CK => CLK, RN => 
                           n2965, Q => REGISTERS_84_8_port, QN => n_1307);
   REGISTERS_reg_84_7_inst : DFFR_X1 port map( D => n9029, CK => CLK, RN => 
                           n2965, Q => REGISTERS_84_7_port, QN => n_1308);
   REGISTERS_reg_84_6_inst : DFFR_X1 port map( D => n9030, CK => CLK, RN => 
                           n2965, Q => REGISTERS_84_6_port, QN => n_1309);
   REGISTERS_reg_84_5_inst : DFFR_X1 port map( D => n9031, CK => CLK, RN => 
                           n2965, Q => REGISTERS_84_5_port, QN => n_1310);
   REGISTERS_reg_84_4_inst : DFFR_X1 port map( D => n9032, CK => CLK, RN => 
                           n2965, Q => REGISTERS_84_4_port, QN => n_1311);
   REGISTERS_reg_84_3_inst : DFFR_X1 port map( D => n9033, CK => CLK, RN => 
                           n2964, Q => REGISTERS_84_3_port, QN => n_1312);
   REGISTERS_reg_84_2_inst : DFFR_X1 port map( D => n9034, CK => CLK, RN => 
                           n2964, Q => REGISTERS_84_2_port, QN => n_1313);
   REGISTERS_reg_84_1_inst : DFFR_X1 port map( D => n9035, CK => CLK, RN => 
                           n2964, Q => REGISTERS_84_1_port, QN => n_1314);
   REGISTERS_reg_84_0_inst : DFFR_X1 port map( D => n9036, CK => CLK, RN => 
                           n2964, Q => REGISTERS_84_0_port, QN => n_1315);
   REGISTERS_reg_83_31_inst : DFFR_X1 port map( D => n8973, CK => CLK, RN => 
                           n2969, Q => REGISTERS_83_31_port, QN => n_1316);
   REGISTERS_reg_83_30_inst : DFFR_X1 port map( D => n8974, CK => CLK, RN => 
                           n2969, Q => REGISTERS_83_30_port, QN => n_1317);
   REGISTERS_reg_83_29_inst : DFFR_X1 port map( D => n8975, CK => CLK, RN => 
                           n2969, Q => REGISTERS_83_29_port, QN => n_1318);
   REGISTERS_reg_83_28_inst : DFFR_X1 port map( D => n8976, CK => CLK, RN => 
                           n2969, Q => REGISTERS_83_28_port, QN => n_1319);
   REGISTERS_reg_83_27_inst : DFFR_X1 port map( D => n8977, CK => CLK, RN => 
                           n2969, Q => REGISTERS_83_27_port, QN => n_1320);
   REGISTERS_reg_83_26_inst : DFFR_X1 port map( D => n8978, CK => CLK, RN => 
                           n2969, Q => REGISTERS_83_26_port, QN => n_1321);
   REGISTERS_reg_83_25_inst : DFFR_X1 port map( D => n8979, CK => CLK, RN => 
                           n2969, Q => REGISTERS_83_25_port, QN => n_1322);
   REGISTERS_reg_83_24_inst : DFFR_X1 port map( D => n8980, CK => CLK, RN => 
                           n2969, Q => REGISTERS_83_24_port, QN => n_1323);
   REGISTERS_reg_83_23_inst : DFFR_X1 port map( D => n8981, CK => CLK, RN => 
                           n2969, Q => REGISTERS_83_23_port, QN => n_1324);
   REGISTERS_reg_83_22_inst : DFFR_X1 port map( D => n8982, CK => CLK, RN => 
                           n2969, Q => REGISTERS_83_22_port, QN => n_1325);
   REGISTERS_reg_83_21_inst : DFFR_X1 port map( D => n8983, CK => CLK, RN => 
                           n2969, Q => REGISTERS_83_21_port, QN => n_1326);
   REGISTERS_reg_83_20_inst : DFFR_X1 port map( D => n8984, CK => CLK, RN => 
                           n2969, Q => REGISTERS_83_20_port, QN => n_1327);
   REGISTERS_reg_83_19_inst : DFFR_X1 port map( D => n8985, CK => CLK, RN => 
                           n2968, Q => REGISTERS_83_19_port, QN => n_1328);
   REGISTERS_reg_83_18_inst : DFFR_X1 port map( D => n8986, CK => CLK, RN => 
                           n2968, Q => REGISTERS_83_18_port, QN => n_1329);
   REGISTERS_reg_83_17_inst : DFFR_X1 port map( D => n8987, CK => CLK, RN => 
                           n2968, Q => REGISTERS_83_17_port, QN => n_1330);
   REGISTERS_reg_83_16_inst : DFFR_X1 port map( D => n8988, CK => CLK, RN => 
                           n2968, Q => REGISTERS_83_16_port, QN => n_1331);
   REGISTERS_reg_83_15_inst : DFFR_X1 port map( D => n8989, CK => CLK, RN => 
                           n2968, Q => REGISTERS_83_15_port, QN => n_1332);
   REGISTERS_reg_83_14_inst : DFFR_X1 port map( D => n8990, CK => CLK, RN => 
                           n2968, Q => REGISTERS_83_14_port, QN => n_1333);
   REGISTERS_reg_83_13_inst : DFFR_X1 port map( D => n8991, CK => CLK, RN => 
                           n2968, Q => REGISTERS_83_13_port, QN => n_1334);
   REGISTERS_reg_83_12_inst : DFFR_X1 port map( D => n8992, CK => CLK, RN => 
                           n2968, Q => REGISTERS_83_12_port, QN => n_1335);
   REGISTERS_reg_83_11_inst : DFFR_X1 port map( D => n8993, CK => CLK, RN => 
                           n2968, Q => REGISTERS_83_11_port, QN => n_1336);
   REGISTERS_reg_83_10_inst : DFFR_X1 port map( D => n8994, CK => CLK, RN => 
                           n2968, Q => REGISTERS_83_10_port, QN => n_1337);
   REGISTERS_reg_83_9_inst : DFFR_X1 port map( D => n8995, CK => CLK, RN => 
                           n2968, Q => REGISTERS_83_9_port, QN => n_1338);
   REGISTERS_reg_83_8_inst : DFFR_X1 port map( D => n8996, CK => CLK, RN => 
                           n2968, Q => REGISTERS_83_8_port, QN => n_1339);
   REGISTERS_reg_83_7_inst : DFFR_X1 port map( D => n8997, CK => CLK, RN => 
                           n2967, Q => REGISTERS_83_7_port, QN => n_1340);
   REGISTERS_reg_83_6_inst : DFFR_X1 port map( D => n8998, CK => CLK, RN => 
                           n2967, Q => REGISTERS_83_6_port, QN => n_1341);
   REGISTERS_reg_83_5_inst : DFFR_X1 port map( D => n8999, CK => CLK, RN => 
                           n2967, Q => REGISTERS_83_5_port, QN => n_1342);
   REGISTERS_reg_83_4_inst : DFFR_X1 port map( D => n9000, CK => CLK, RN => 
                           n2967, Q => REGISTERS_83_4_port, QN => n_1343);
   REGISTERS_reg_83_3_inst : DFFR_X1 port map( D => n9001, CK => CLK, RN => 
                           n2967, Q => REGISTERS_83_3_port, QN => n_1344);
   REGISTERS_reg_83_2_inst : DFFR_X1 port map( D => n9002, CK => CLK, RN => 
                           n2967, Q => REGISTERS_83_2_port, QN => n_1345);
   REGISTERS_reg_83_1_inst : DFFR_X1 port map( D => n9003, CK => CLK, RN => 
                           n2967, Q => REGISTERS_83_1_port, QN => n_1346);
   REGISTERS_reg_83_0_inst : DFFR_X1 port map( D => n9004, CK => CLK, RN => 
                           n2967, Q => REGISTERS_83_0_port, QN => n_1347);
   REGISTERS_reg_82_31_inst : DFFR_X1 port map( D => n8941, CK => CLK, RN => 
                           n2972, Q => REGISTERS_82_31_port, QN => n_1348);
   REGISTERS_reg_82_30_inst : DFFR_X1 port map( D => n8942, CK => CLK, RN => 
                           n2972, Q => REGISTERS_82_30_port, QN => n_1349);
   REGISTERS_reg_82_29_inst : DFFR_X1 port map( D => n8943, CK => CLK, RN => 
                           n2972, Q => REGISTERS_82_29_port, QN => n_1350);
   REGISTERS_reg_82_28_inst : DFFR_X1 port map( D => n8944, CK => CLK, RN => 
                           n2972, Q => REGISTERS_82_28_port, QN => n_1351);
   REGISTERS_reg_82_27_inst : DFFR_X1 port map( D => n8945, CK => CLK, RN => 
                           n2972, Q => REGISTERS_82_27_port, QN => n_1352);
   REGISTERS_reg_82_26_inst : DFFR_X1 port map( D => n8946, CK => CLK, RN => 
                           n2972, Q => REGISTERS_82_26_port, QN => n_1353);
   REGISTERS_reg_82_25_inst : DFFR_X1 port map( D => n8947, CK => CLK, RN => 
                           n2972, Q => REGISTERS_82_25_port, QN => n_1354);
   REGISTERS_reg_82_24_inst : DFFR_X1 port map( D => n8948, CK => CLK, RN => 
                           n2972, Q => REGISTERS_82_24_port, QN => n_1355);
   REGISTERS_reg_82_23_inst : DFFR_X1 port map( D => n8949, CK => CLK, RN => 
                           n2971, Q => REGISTERS_82_23_port, QN => n_1356);
   REGISTERS_reg_82_22_inst : DFFR_X1 port map( D => n8950, CK => CLK, RN => 
                           n2971, Q => REGISTERS_82_22_port, QN => n_1357);
   REGISTERS_reg_82_21_inst : DFFR_X1 port map( D => n8951, CK => CLK, RN => 
                           n2971, Q => REGISTERS_82_21_port, QN => n_1358);
   REGISTERS_reg_82_20_inst : DFFR_X1 port map( D => n8952, CK => CLK, RN => 
                           n2971, Q => REGISTERS_82_20_port, QN => n_1359);
   REGISTERS_reg_82_19_inst : DFFR_X1 port map( D => n8953, CK => CLK, RN => 
                           n2971, Q => REGISTERS_82_19_port, QN => n_1360);
   REGISTERS_reg_82_18_inst : DFFR_X1 port map( D => n8954, CK => CLK, RN => 
                           n2971, Q => REGISTERS_82_18_port, QN => n_1361);
   REGISTERS_reg_82_17_inst : DFFR_X1 port map( D => n8955, CK => CLK, RN => 
                           n2971, Q => REGISTERS_82_17_port, QN => n_1362);
   REGISTERS_reg_82_16_inst : DFFR_X1 port map( D => n8956, CK => CLK, RN => 
                           n2971, Q => REGISTERS_82_16_port, QN => n_1363);
   REGISTERS_reg_82_15_inst : DFFR_X1 port map( D => n8957, CK => CLK, RN => 
                           n2971, Q => REGISTERS_82_15_port, QN => n_1364);
   REGISTERS_reg_82_14_inst : DFFR_X1 port map( D => n8958, CK => CLK, RN => 
                           n2971, Q => REGISTERS_82_14_port, QN => n_1365);
   REGISTERS_reg_82_13_inst : DFFR_X1 port map( D => n8959, CK => CLK, RN => 
                           n2971, Q => REGISTERS_82_13_port, QN => n_1366);
   REGISTERS_reg_82_12_inst : DFFR_X1 port map( D => n8960, CK => CLK, RN => 
                           n2971, Q => REGISTERS_82_12_port, QN => n_1367);
   REGISTERS_reg_82_11_inst : DFFR_X1 port map( D => n8961, CK => CLK, RN => 
                           n2970, Q => REGISTERS_82_11_port, QN => n_1368);
   REGISTERS_reg_82_10_inst : DFFR_X1 port map( D => n8962, CK => CLK, RN => 
                           n2970, Q => REGISTERS_82_10_port, QN => n_1369);
   REGISTERS_reg_82_9_inst : DFFR_X1 port map( D => n8963, CK => CLK, RN => 
                           n2970, Q => REGISTERS_82_9_port, QN => n_1370);
   REGISTERS_reg_82_8_inst : DFFR_X1 port map( D => n8964, CK => CLK, RN => 
                           n2970, Q => REGISTERS_82_8_port, QN => n_1371);
   REGISTERS_reg_82_7_inst : DFFR_X1 port map( D => n8965, CK => CLK, RN => 
                           n2970, Q => REGISTERS_82_7_port, QN => n_1372);
   REGISTERS_reg_82_6_inst : DFFR_X1 port map( D => n8966, CK => CLK, RN => 
                           n2970, Q => REGISTERS_82_6_port, QN => n_1373);
   REGISTERS_reg_82_5_inst : DFFR_X1 port map( D => n8967, CK => CLK, RN => 
                           n2970, Q => REGISTERS_82_5_port, QN => n_1374);
   REGISTERS_reg_82_4_inst : DFFR_X1 port map( D => n8968, CK => CLK, RN => 
                           n2970, Q => REGISTERS_82_4_port, QN => n_1375);
   REGISTERS_reg_82_3_inst : DFFR_X1 port map( D => n8969, CK => CLK, RN => 
                           n2970, Q => REGISTERS_82_3_port, QN => n_1376);
   REGISTERS_reg_82_2_inst : DFFR_X1 port map( D => n8970, CK => CLK, RN => 
                           n2970, Q => REGISTERS_82_2_port, QN => n_1377);
   REGISTERS_reg_82_1_inst : DFFR_X1 port map( D => n8971, CK => CLK, RN => 
                           n2970, Q => REGISTERS_82_1_port, QN => n_1378);
   REGISTERS_reg_82_0_inst : DFFR_X1 port map( D => n8972, CK => CLK, RN => 
                           n2970, Q => REGISTERS_82_0_port, QN => n_1379);
   REGISTERS_reg_78_31_inst : DFFR_X1 port map( D => n8813, CK => CLK, RN => 
                           n2983, Q => REGISTERS_78_31_port, QN => n_1380);
   REGISTERS_reg_78_30_inst : DFFR_X1 port map( D => n8814, CK => CLK, RN => 
                           n2983, Q => REGISTERS_78_30_port, QN => n_1381);
   REGISTERS_reg_78_29_inst : DFFR_X1 port map( D => n8815, CK => CLK, RN => 
                           n2983, Q => REGISTERS_78_29_port, QN => n_1382);
   REGISTERS_reg_78_28_inst : DFFR_X1 port map( D => n8816, CK => CLK, RN => 
                           n2983, Q => REGISTERS_78_28_port, QN => n_1383);
   REGISTERS_reg_78_27_inst : DFFR_X1 port map( D => n8817, CK => CLK, RN => 
                           n2982, Q => REGISTERS_78_27_port, QN => n_1384);
   REGISTERS_reg_78_26_inst : DFFR_X1 port map( D => n8818, CK => CLK, RN => 
                           n2982, Q => REGISTERS_78_26_port, QN => n_1385);
   REGISTERS_reg_78_25_inst : DFFR_X1 port map( D => n8819, CK => CLK, RN => 
                           n2982, Q => REGISTERS_78_25_port, QN => n_1386);
   REGISTERS_reg_78_24_inst : DFFR_X1 port map( D => n8820, CK => CLK, RN => 
                           n2982, Q => REGISTERS_78_24_port, QN => n_1387);
   REGISTERS_reg_78_23_inst : DFFR_X1 port map( D => n8821, CK => CLK, RN => 
                           n2982, Q => REGISTERS_78_23_port, QN => n_1388);
   REGISTERS_reg_78_22_inst : DFFR_X1 port map( D => n8822, CK => CLK, RN => 
                           n2982, Q => REGISTERS_78_22_port, QN => n_1389);
   REGISTERS_reg_78_21_inst : DFFR_X1 port map( D => n8823, CK => CLK, RN => 
                           n2982, Q => REGISTERS_78_21_port, QN => n_1390);
   REGISTERS_reg_78_20_inst : DFFR_X1 port map( D => n8824, CK => CLK, RN => 
                           n2982, Q => REGISTERS_78_20_port, QN => n_1391);
   REGISTERS_reg_78_19_inst : DFFR_X1 port map( D => n8825, CK => CLK, RN => 
                           n2982, Q => REGISTERS_78_19_port, QN => n_1392);
   REGISTERS_reg_78_18_inst : DFFR_X1 port map( D => n8826, CK => CLK, RN => 
                           n2982, Q => REGISTERS_78_18_port, QN => n_1393);
   REGISTERS_reg_78_17_inst : DFFR_X1 port map( D => n8827, CK => CLK, RN => 
                           n2982, Q => REGISTERS_78_17_port, QN => n_1394);
   REGISTERS_reg_78_16_inst : DFFR_X1 port map( D => n8828, CK => CLK, RN => 
                           n2982, Q => REGISTERS_78_16_port, QN => n_1395);
   REGISTERS_reg_78_15_inst : DFFR_X1 port map( D => n8829, CK => CLK, RN => 
                           n2981, Q => REGISTERS_78_15_port, QN => n_1396);
   REGISTERS_reg_78_14_inst : DFFR_X1 port map( D => n8830, CK => CLK, RN => 
                           n2981, Q => REGISTERS_78_14_port, QN => n_1397);
   REGISTERS_reg_78_13_inst : DFFR_X1 port map( D => n8831, CK => CLK, RN => 
                           n2981, Q => REGISTERS_78_13_port, QN => n_1398);
   REGISTERS_reg_78_12_inst : DFFR_X1 port map( D => n8832, CK => CLK, RN => 
                           n2981, Q => REGISTERS_78_12_port, QN => n_1399);
   REGISTERS_reg_78_11_inst : DFFR_X1 port map( D => n8833_port, CK => CLK, RN 
                           => n2981, Q => REGISTERS_78_11_port, QN => n_1400);
   REGISTERS_reg_78_10_inst : DFFR_X1 port map( D => n8834_port, CK => CLK, RN 
                           => n2981, Q => REGISTERS_78_10_port, QN => n_1401);
   REGISTERS_reg_78_9_inst : DFFR_X1 port map( D => n8835, CK => CLK, RN => 
                           n2981, Q => REGISTERS_78_9_port, QN => n_1402);
   REGISTERS_reg_78_8_inst : DFFR_X1 port map( D => n8836, CK => CLK, RN => 
                           n2981, Q => REGISTERS_78_8_port, QN => n_1403);
   REGISTERS_reg_78_7_inst : DFFR_X1 port map( D => n8837, CK => CLK, RN => 
                           n2981, Q => REGISTERS_78_7_port, QN => n_1404);
   REGISTERS_reg_78_6_inst : DFFR_X1 port map( D => n8838, CK => CLK, RN => 
                           n2981, Q => REGISTERS_78_6_port, QN => n_1405);
   REGISTERS_reg_78_5_inst : DFFR_X1 port map( D => n8839, CK => CLK, RN => 
                           n2981, Q => REGISTERS_78_5_port, QN => n_1406);
   REGISTERS_reg_78_4_inst : DFFR_X1 port map( D => n8840, CK => CLK, RN => 
                           n2981, Q => REGISTERS_78_4_port, QN => n_1407);
   REGISTERS_reg_78_3_inst : DFFR_X1 port map( D => n8841, CK => CLK, RN => 
                           n2980, Q => REGISTERS_78_3_port, QN => n_1408);
   REGISTERS_reg_78_2_inst : DFFR_X1 port map( D => n8842, CK => CLK, RN => 
                           n2980, Q => REGISTERS_78_2_port, QN => n_1409);
   REGISTERS_reg_78_1_inst : DFFR_X1 port map( D => n8843, CK => CLK, RN => 
                           n2980, Q => REGISTERS_78_1_port, QN => n_1410);
   REGISTERS_reg_78_0_inst : DFFR_X1 port map( D => n8844, CK => CLK, RN => 
                           n2980, Q => REGISTERS_78_0_port, QN => n_1411);
   REGISTERS_reg_77_31_inst : DFFR_X1 port map( D => n8781, CK => CLK, RN => 
                           n2985, Q => REGISTERS_77_31_port, QN => n_1412);
   REGISTERS_reg_77_30_inst : DFFR_X1 port map( D => n8782, CK => CLK, RN => 
                           n2985, Q => REGISTERS_77_30_port, QN => n_1413);
   REGISTERS_reg_77_29_inst : DFFR_X1 port map( D => n8783, CK => CLK, RN => 
                           n2985, Q => REGISTERS_77_29_port, QN => n_1414);
   REGISTERS_reg_77_28_inst : DFFR_X1 port map( D => n8784, CK => CLK, RN => 
                           n2985, Q => REGISTERS_77_28_port, QN => n_1415);
   REGISTERS_reg_77_27_inst : DFFR_X1 port map( D => n8785, CK => CLK, RN => 
                           n2985, Q => REGISTERS_77_27_port, QN => n_1416);
   REGISTERS_reg_77_26_inst : DFFR_X1 port map( D => n8786, CK => CLK, RN => 
                           n2985, Q => REGISTERS_77_26_port, QN => n_1417);
   REGISTERS_reg_77_25_inst : DFFR_X1 port map( D => n8787_port, CK => CLK, RN 
                           => n2985, Q => REGISTERS_77_25_port, QN => n_1418);
   REGISTERS_reg_77_24_inst : DFFR_X1 port map( D => n8788_port, CK => CLK, RN 
                           => n2985, Q => REGISTERS_77_24_port, QN => n_1419);
   REGISTERS_reg_77_23_inst : DFFR_X1 port map( D => n8789_port, CK => CLK, RN 
                           => n2985, Q => REGISTERS_77_23_port, QN => n_1420);
   REGISTERS_reg_77_22_inst : DFFR_X1 port map( D => n8790_port, CK => CLK, RN 
                           => n2985, Q => REGISTERS_77_22_port, QN => n_1421);
   REGISTERS_reg_77_21_inst : DFFR_X1 port map( D => n8791_port, CK => CLK, RN 
                           => n2985, Q => REGISTERS_77_21_port, QN => n_1422);
   REGISTERS_reg_77_20_inst : DFFR_X1 port map( D => n8792, CK => CLK, RN => 
                           n2985, Q => REGISTERS_77_20_port, QN => n_1423);
   REGISTERS_reg_77_19_inst : DFFR_X1 port map( D => n8793, CK => CLK, RN => 
                           n2984, Q => REGISTERS_77_19_port, QN => n_1424);
   REGISTERS_reg_77_18_inst : DFFR_X1 port map( D => n8794, CK => CLK, RN => 
                           n2984, Q => REGISTERS_77_18_port, QN => n_1425);
   REGISTERS_reg_77_17_inst : DFFR_X1 port map( D => n8795, CK => CLK, RN => 
                           n2984, Q => REGISTERS_77_17_port, QN => n_1426);
   REGISTERS_reg_77_16_inst : DFFR_X1 port map( D => n8796, CK => CLK, RN => 
                           n2984, Q => REGISTERS_77_16_port, QN => n_1427);
   REGISTERS_reg_77_15_inst : DFFR_X1 port map( D => n8797, CK => CLK, RN => 
                           n2984, Q => REGISTERS_77_15_port, QN => n_1428);
   REGISTERS_reg_77_14_inst : DFFR_X1 port map( D => n8798, CK => CLK, RN => 
                           n2984, Q => REGISTERS_77_14_port, QN => n_1429);
   REGISTERS_reg_77_13_inst : DFFR_X1 port map( D => n8799, CK => CLK, RN => 
                           n2984, Q => REGISTERS_77_13_port, QN => n_1430);
   REGISTERS_reg_77_12_inst : DFFR_X1 port map( D => n8800, CK => CLK, RN => 
                           n2984, Q => REGISTERS_77_12_port, QN => n_1431);
   REGISTERS_reg_77_11_inst : DFFR_X1 port map( D => n8801, CK => CLK, RN => 
                           n2984, Q => REGISTERS_77_11_port, QN => n_1432);
   REGISTERS_reg_77_10_inst : DFFR_X1 port map( D => n8802, CK => CLK, RN => 
                           n2984, Q => REGISTERS_77_10_port, QN => n_1433);
   REGISTERS_reg_77_9_inst : DFFR_X1 port map( D => n8803, CK => CLK, RN => 
                           n2984, Q => REGISTERS_77_9_port, QN => n_1434);
   REGISTERS_reg_77_8_inst : DFFR_X1 port map( D => n8804, CK => CLK, RN => 
                           n2984, Q => REGISTERS_77_8_port, QN => n_1435);
   REGISTERS_reg_77_7_inst : DFFR_X1 port map( D => n8805, CK => CLK, RN => 
                           n2983, Q => REGISTERS_77_7_port, QN => n_1436);
   REGISTERS_reg_77_6_inst : DFFR_X1 port map( D => n8806, CK => CLK, RN => 
                           n2983, Q => REGISTERS_77_6_port, QN => n_1437);
   REGISTERS_reg_77_5_inst : DFFR_X1 port map( D => n8807, CK => CLK, RN => 
                           n2983, Q => REGISTERS_77_5_port, QN => n_1438);
   REGISTERS_reg_77_4_inst : DFFR_X1 port map( D => n8808, CK => CLK, RN => 
                           n2983, Q => REGISTERS_77_4_port, QN => n_1439);
   REGISTERS_reg_77_3_inst : DFFR_X1 port map( D => n8809, CK => CLK, RN => 
                           n2983, Q => REGISTERS_77_3_port, QN => n_1440);
   REGISTERS_reg_77_2_inst : DFFR_X1 port map( D => n8810, CK => CLK, RN => 
                           n2983, Q => REGISTERS_77_2_port, QN => n_1441);
   REGISTERS_reg_77_1_inst : DFFR_X1 port map( D => n8811, CK => CLK, RN => 
                           n2983, Q => REGISTERS_77_1_port, QN => n_1442);
   REGISTERS_reg_77_0_inst : DFFR_X1 port map( D => n8812, CK => CLK, RN => 
                           n2983, Q => REGISTERS_77_0_port, QN => n_1443);
   REGISTERS_reg_54_31_inst : DFFR_X1 port map( D => n8045, CK => CLK, RN => 
                           n3061, Q => REGISTERS_54_31_port, QN => n_1444);
   REGISTERS_reg_54_30_inst : DFFR_X1 port map( D => n8046, CK => CLK, RN => 
                           n3061, Q => REGISTERS_54_30_port, QN => n_1445);
   REGISTERS_reg_54_29_inst : DFFR_X1 port map( D => n8047, CK => CLK, RN => 
                           n3061, Q => REGISTERS_54_29_port, QN => n_1446);
   REGISTERS_reg_54_28_inst : DFFR_X1 port map( D => n8048, CK => CLK, RN => 
                           n3061, Q => REGISTERS_54_28_port, QN => n_1447);
   REGISTERS_reg_54_27_inst : DFFR_X1 port map( D => n8049, CK => CLK, RN => 
                           n3059, Q => REGISTERS_54_27_port, QN => n_1448);
   REGISTERS_reg_54_26_inst : DFFR_X1 port map( D => n8050, CK => CLK, RN => 
                           n3059, Q => REGISTERS_54_26_port, QN => n_1449);
   REGISTERS_reg_54_25_inst : DFFR_X1 port map( D => n8051, CK => CLK, RN => 
                           n3059, Q => REGISTERS_54_25_port, QN => n_1450);
   REGISTERS_reg_54_24_inst : DFFR_X1 port map( D => n8052, CK => CLK, RN => 
                           n3059, Q => REGISTERS_54_24_port, QN => n_1451);
   REGISTERS_reg_54_23_inst : DFFR_X1 port map( D => n8053, CK => CLK, RN => 
                           n3059, Q => REGISTERS_54_23_port, QN => n_1452);
   REGISTERS_reg_54_22_inst : DFFR_X1 port map( D => n8054, CK => CLK, RN => 
                           n3059, Q => REGISTERS_54_22_port, QN => n_1453);
   REGISTERS_reg_54_21_inst : DFFR_X1 port map( D => n8055, CK => CLK, RN => 
                           n3059, Q => REGISTERS_54_21_port, QN => n_1454);
   REGISTERS_reg_54_20_inst : DFFR_X1 port map( D => n8056, CK => CLK, RN => 
                           n3059, Q => REGISTERS_54_20_port, QN => n_1455);
   REGISTERS_reg_54_19_inst : DFFR_X1 port map( D => n8057, CK => CLK, RN => 
                           n3059, Q => REGISTERS_54_19_port, QN => n_1456);
   REGISTERS_reg_54_18_inst : DFFR_X1 port map( D => n8058, CK => CLK, RN => 
                           n3059, Q => REGISTERS_54_18_port, QN => n_1457);
   REGISTERS_reg_54_17_inst : DFFR_X1 port map( D => n8059, CK => CLK, RN => 
                           n3059, Q => REGISTERS_54_17_port, QN => n_1458);
   REGISTERS_reg_54_16_inst : DFFR_X1 port map( D => n8060, CK => CLK, RN => 
                           n3059, Q => REGISTERS_54_16_port, QN => n_1459);
   REGISTERS_reg_54_15_inst : DFFR_X1 port map( D => n8061, CK => CLK, RN => 
                           n3057, Q => REGISTERS_54_15_port, QN => n_1460);
   REGISTERS_reg_54_14_inst : DFFR_X1 port map( D => n8062, CK => CLK, RN => 
                           n3057, Q => REGISTERS_54_14_port, QN => n_1461);
   REGISTERS_reg_54_13_inst : DFFR_X1 port map( D => n8063, CK => CLK, RN => 
                           n3057, Q => REGISTERS_54_13_port, QN => n_1462);
   REGISTERS_reg_54_12_inst : DFFR_X1 port map( D => n8064, CK => CLK, RN => 
                           n3057, Q => REGISTERS_54_12_port, QN => n_1463);
   REGISTERS_reg_54_11_inst : DFFR_X1 port map( D => n8065, CK => CLK, RN => 
                           n3057, Q => REGISTERS_54_11_port, QN => n_1464);
   REGISTERS_reg_54_10_inst : DFFR_X1 port map( D => n8066, CK => CLK, RN => 
                           n3057, Q => REGISTERS_54_10_port, QN => n_1465);
   REGISTERS_reg_54_9_inst : DFFR_X1 port map( D => n8067, CK => CLK, RN => 
                           n3057, Q => REGISTERS_54_9_port, QN => n_1466);
   REGISTERS_reg_54_8_inst : DFFR_X1 port map( D => n8068, CK => CLK, RN => 
                           n3057, Q => REGISTERS_54_8_port, QN => n_1467);
   REGISTERS_reg_54_7_inst : DFFR_X1 port map( D => n8069, CK => CLK, RN => 
                           n3057, Q => REGISTERS_54_7_port, QN => n_1468);
   REGISTERS_reg_54_6_inst : DFFR_X1 port map( D => n8070, CK => CLK, RN => 
                           n3057, Q => REGISTERS_54_6_port, QN => n_1469);
   REGISTERS_reg_54_5_inst : DFFR_X1 port map( D => n8071, CK => CLK, RN => 
                           n3057, Q => REGISTERS_54_5_port, QN => n_1470);
   REGISTERS_reg_54_4_inst : DFFR_X1 port map( D => n8072, CK => CLK, RN => 
                           n3057, Q => REGISTERS_54_4_port, QN => n_1471);
   REGISTERS_reg_54_3_inst : DFFR_X1 port map( D => n8073, CK => CLK, RN => 
                           n3056, Q => REGISTERS_54_3_port, QN => n_1472);
   REGISTERS_reg_54_2_inst : DFFR_X1 port map( D => n8074, CK => CLK, RN => 
                           n3056, Q => REGISTERS_54_2_port, QN => n_1473);
   REGISTERS_reg_54_1_inst : DFFR_X1 port map( D => n8075, CK => CLK, RN => 
                           n3056, Q => REGISTERS_54_1_port, QN => n_1474);
   REGISTERS_reg_54_0_inst : DFFR_X1 port map( D => n8076, CK => CLK, RN => 
                           n3056, Q => REGISTERS_54_0_port, QN => n_1475);
   REGISTERS_reg_53_31_inst : DFFR_X1 port map( D => n8013, CK => CLK, RN => 
                           n3064, Q => REGISTERS_53_31_port, QN => n_1476);
   REGISTERS_reg_53_30_inst : DFFR_X1 port map( D => n8014, CK => CLK, RN => 
                           n3064, Q => REGISTERS_53_30_port, QN => n_1477);
   REGISTERS_reg_53_29_inst : DFFR_X1 port map( D => n8015, CK => CLK, RN => 
                           n3064, Q => REGISTERS_53_29_port, QN => n_1478);
   REGISTERS_reg_53_28_inst : DFFR_X1 port map( D => n8016, CK => CLK, RN => 
                           n3064, Q => REGISTERS_53_28_port, QN => n_1479);
   REGISTERS_reg_53_27_inst : DFFR_X1 port map( D => n8017, CK => CLK, RN => 
                           n3064, Q => REGISTERS_53_27_port, QN => n_1480);
   REGISTERS_reg_53_26_inst : DFFR_X1 port map( D => n8018, CK => CLK, RN => 
                           n3064, Q => REGISTERS_53_26_port, QN => n_1481);
   REGISTERS_reg_53_25_inst : DFFR_X1 port map( D => n8019, CK => CLK, RN => 
                           n3064, Q => REGISTERS_53_25_port, QN => n_1482);
   REGISTERS_reg_53_24_inst : DFFR_X1 port map( D => n8020, CK => CLK, RN => 
                           n3064, Q => REGISTERS_53_24_port, QN => n_1483);
   REGISTERS_reg_53_23_inst : DFFR_X1 port map( D => n8021, CK => CLK, RN => 
                           n3064, Q => REGISTERS_53_23_port, QN => n_1484);
   REGISTERS_reg_53_22_inst : DFFR_X1 port map( D => n8022, CK => CLK, RN => 
                           n3064, Q => REGISTERS_53_22_port, QN => n_1485);
   REGISTERS_reg_53_21_inst : DFFR_X1 port map( D => n8023, CK => CLK, RN => 
                           n3064, Q => REGISTERS_53_21_port, QN => n_1486);
   REGISTERS_reg_53_20_inst : DFFR_X1 port map( D => n8024, CK => CLK, RN => 
                           n3064, Q => REGISTERS_53_20_port, QN => n_1487);
   REGISTERS_reg_53_19_inst : DFFR_X1 port map( D => n8025, CK => CLK, RN => 
                           n3062, Q => REGISTERS_53_19_port, QN => n_1488);
   REGISTERS_reg_53_18_inst : DFFR_X1 port map( D => n8026, CK => CLK, RN => 
                           n3062, Q => REGISTERS_53_18_port, QN => n_1489);
   REGISTERS_reg_53_17_inst : DFFR_X1 port map( D => n8027, CK => CLK, RN => 
                           n3062, Q => REGISTERS_53_17_port, QN => n_1490);
   REGISTERS_reg_53_16_inst : DFFR_X1 port map( D => n8028, CK => CLK, RN => 
                           n3062, Q => REGISTERS_53_16_port, QN => n_1491);
   REGISTERS_reg_53_15_inst : DFFR_X1 port map( D => n8029, CK => CLK, RN => 
                           n3062, Q => REGISTERS_53_15_port, QN => n_1492);
   REGISTERS_reg_53_14_inst : DFFR_X1 port map( D => n8030, CK => CLK, RN => 
                           n3062, Q => REGISTERS_53_14_port, QN => n_1493);
   REGISTERS_reg_53_13_inst : DFFR_X1 port map( D => n8031, CK => CLK, RN => 
                           n3062, Q => REGISTERS_53_13_port, QN => n_1494);
   REGISTERS_reg_53_12_inst : DFFR_X1 port map( D => n8032, CK => CLK, RN => 
                           n3062, Q => REGISTERS_53_12_port, QN => n_1495);
   REGISTERS_reg_53_11_inst : DFFR_X1 port map( D => n8033, CK => CLK, RN => 
                           n3062, Q => REGISTERS_53_11_port, QN => n_1496);
   REGISTERS_reg_53_10_inst : DFFR_X1 port map( D => n8034, CK => CLK, RN => 
                           n3062, Q => REGISTERS_53_10_port, QN => n_1497);
   REGISTERS_reg_53_9_inst : DFFR_X1 port map( D => n8035, CK => CLK, RN => 
                           n3062, Q => REGISTERS_53_9_port, QN => n_1498);
   REGISTERS_reg_53_8_inst : DFFR_X1 port map( D => n8036, CK => CLK, RN => 
                           n3062, Q => REGISTERS_53_8_port, QN => n_1499);
   REGISTERS_reg_53_7_inst : DFFR_X1 port map( D => n8037, CK => CLK, RN => 
                           n3061, Q => REGISTERS_53_7_port, QN => n_1500);
   REGISTERS_reg_53_6_inst : DFFR_X1 port map( D => n8038, CK => CLK, RN => 
                           n3061, Q => REGISTERS_53_6_port, QN => n_1501);
   REGISTERS_reg_53_5_inst : DFFR_X1 port map( D => n8039, CK => CLK, RN => 
                           n3061, Q => REGISTERS_53_5_port, QN => n_1502);
   REGISTERS_reg_53_4_inst : DFFR_X1 port map( D => n8040, CK => CLK, RN => 
                           n3061, Q => REGISTERS_53_4_port, QN => n_1503);
   REGISTERS_reg_53_3_inst : DFFR_X1 port map( D => n8041, CK => CLK, RN => 
                           n3061, Q => REGISTERS_53_3_port, QN => n_1504);
   REGISTERS_reg_53_2_inst : DFFR_X1 port map( D => n8042, CK => CLK, RN => 
                           n3061, Q => REGISTERS_53_2_port, QN => n_1505);
   REGISTERS_reg_53_1_inst : DFFR_X1 port map( D => n8043, CK => CLK, RN => 
                           n3061, Q => REGISTERS_53_1_port, QN => n_1506);
   REGISTERS_reg_53_0_inst : DFFR_X1 port map( D => n8044, CK => CLK, RN => 
                           n3061, Q => REGISTERS_53_0_port, QN => n_1507);
   REGISTERS_reg_52_31_inst : DFFR_X1 port map( D => n7981, CK => CLK, RN => 
                           n3069, Q => REGISTERS_52_31_port, QN => n_1508);
   REGISTERS_reg_52_30_inst : DFFR_X1 port map( D => n7982, CK => CLK, RN => 
                           n3069, Q => REGISTERS_52_30_port, QN => n_1509);
   REGISTERS_reg_52_29_inst : DFFR_X1 port map( D => n7983, CK => CLK, RN => 
                           n3069, Q => REGISTERS_52_29_port, QN => n_1510);
   REGISTERS_reg_52_28_inst : DFFR_X1 port map( D => n7984, CK => CLK, RN => 
                           n3069, Q => REGISTERS_52_28_port, QN => n_1511);
   REGISTERS_reg_52_27_inst : DFFR_X1 port map( D => n7985, CK => CLK, RN => 
                           n3069, Q => REGISTERS_52_27_port, QN => n_1512);
   REGISTERS_reg_52_26_inst : DFFR_X1 port map( D => n7986, CK => CLK, RN => 
                           n3069, Q => REGISTERS_52_26_port, QN => n_1513);
   REGISTERS_reg_52_25_inst : DFFR_X1 port map( D => n7987, CK => CLK, RN => 
                           n3069, Q => REGISTERS_52_25_port, QN => n_1514);
   REGISTERS_reg_52_24_inst : DFFR_X1 port map( D => n7988, CK => CLK, RN => 
                           n3069, Q => REGISTERS_52_24_port, QN => n_1515);
   REGISTERS_reg_52_23_inst : DFFR_X1 port map( D => n7989, CK => CLK, RN => 
                           n3067, Q => REGISTERS_52_23_port, QN => n_1516);
   REGISTERS_reg_52_22_inst : DFFR_X1 port map( D => n7990, CK => CLK, RN => 
                           n3067, Q => REGISTERS_52_22_port, QN => n_1517);
   REGISTERS_reg_52_21_inst : DFFR_X1 port map( D => n7991, CK => CLK, RN => 
                           n3067, Q => REGISTERS_52_21_port, QN => n_1518);
   REGISTERS_reg_52_20_inst : DFFR_X1 port map( D => n7992, CK => CLK, RN => 
                           n3067, Q => REGISTERS_52_20_port, QN => n_1519);
   REGISTERS_reg_52_19_inst : DFFR_X1 port map( D => n7993, CK => CLK, RN => 
                           n3067, Q => REGISTERS_52_19_port, QN => n_1520);
   REGISTERS_reg_52_18_inst : DFFR_X1 port map( D => n7994, CK => CLK, RN => 
                           n3067, Q => REGISTERS_52_18_port, QN => n_1521);
   REGISTERS_reg_52_17_inst : DFFR_X1 port map( D => n7995, CK => CLK, RN => 
                           n3067, Q => REGISTERS_52_17_port, QN => n_1522);
   REGISTERS_reg_52_16_inst : DFFR_X1 port map( D => n7996, CK => CLK, RN => 
                           n3067, Q => REGISTERS_52_16_port, QN => n_1523);
   REGISTERS_reg_52_15_inst : DFFR_X1 port map( D => n7997, CK => CLK, RN => 
                           n3067, Q => REGISTERS_52_15_port, QN => n_1524);
   REGISTERS_reg_52_14_inst : DFFR_X1 port map( D => n7998, CK => CLK, RN => 
                           n3067, Q => REGISTERS_52_14_port, QN => n_1525);
   REGISTERS_reg_52_13_inst : DFFR_X1 port map( D => n7999, CK => CLK, RN => 
                           n3067, Q => REGISTERS_52_13_port, QN => n_1526);
   REGISTERS_reg_52_12_inst : DFFR_X1 port map( D => n8000, CK => CLK, RN => 
                           n3067, Q => REGISTERS_52_12_port, QN => n_1527);
   REGISTERS_reg_52_11_inst : DFFR_X1 port map( D => n8001, CK => CLK, RN => 
                           n3066, Q => REGISTERS_52_11_port, QN => n_1528);
   REGISTERS_reg_52_10_inst : DFFR_X1 port map( D => n8002, CK => CLK, RN => 
                           n3066, Q => REGISTERS_52_10_port, QN => n_1529);
   REGISTERS_reg_52_9_inst : DFFR_X1 port map( D => n8003, CK => CLK, RN => 
                           n3066, Q => REGISTERS_52_9_port, QN => n_1530);
   REGISTERS_reg_52_8_inst : DFFR_X1 port map( D => n8004, CK => CLK, RN => 
                           n3066, Q => REGISTERS_52_8_port, QN => n_1531);
   REGISTERS_reg_52_7_inst : DFFR_X1 port map( D => n8005, CK => CLK, RN => 
                           n3066, Q => REGISTERS_52_7_port, QN => n_1532);
   REGISTERS_reg_52_6_inst : DFFR_X1 port map( D => n8006, CK => CLK, RN => 
                           n3066, Q => REGISTERS_52_6_port, QN => n_1533);
   REGISTERS_reg_52_5_inst : DFFR_X1 port map( D => n8007, CK => CLK, RN => 
                           n3066, Q => REGISTERS_52_5_port, QN => n_1534);
   REGISTERS_reg_52_4_inst : DFFR_X1 port map( D => n8008, CK => CLK, RN => 
                           n3066, Q => REGISTERS_52_4_port, QN => n_1535);
   REGISTERS_reg_52_3_inst : DFFR_X1 port map( D => n8009, CK => CLK, RN => 
                           n3066, Q => REGISTERS_52_3_port, QN => n_1536);
   REGISTERS_reg_52_2_inst : DFFR_X1 port map( D => n8010, CK => CLK, RN => 
                           n3066, Q => REGISTERS_52_2_port, QN => n_1537);
   REGISTERS_reg_52_1_inst : DFFR_X1 port map( D => n8011, CK => CLK, RN => 
                           n3066, Q => REGISTERS_52_1_port, QN => n_1538);
   REGISTERS_reg_52_0_inst : DFFR_X1 port map( D => n8012, CK => CLK, RN => 
                           n3066, Q => REGISTERS_52_0_port, QN => n_1539);
   REGISTERS_reg_51_31_inst : DFFR_X1 port map( D => n7949, CK => CLK, RN => 
                           n3074, Q => REGISTERS_51_31_port, QN => n_1540);
   REGISTERS_reg_51_30_inst : DFFR_X1 port map( D => n7950, CK => CLK, RN => 
                           n3074, Q => REGISTERS_51_30_port, QN => n_1541);
   REGISTERS_reg_51_29_inst : DFFR_X1 port map( D => n7951, CK => CLK, RN => 
                           n3074, Q => REGISTERS_51_29_port, QN => n_1542);
   REGISTERS_reg_51_28_inst : DFFR_X1 port map( D => n7952, CK => CLK, RN => 
                           n3074, Q => REGISTERS_51_28_port, QN => n_1543);
   REGISTERS_reg_51_27_inst : DFFR_X1 port map( D => n7953, CK => CLK, RN => 
                           n3072, Q => REGISTERS_51_27_port, QN => n_1544);
   REGISTERS_reg_51_26_inst : DFFR_X1 port map( D => n7954, CK => CLK, RN => 
                           n3072, Q => REGISTERS_51_26_port, QN => n_1545);
   REGISTERS_reg_51_25_inst : DFFR_X1 port map( D => n7955, CK => CLK, RN => 
                           n3072, Q => REGISTERS_51_25_port, QN => n_1546);
   REGISTERS_reg_51_24_inst : DFFR_X1 port map( D => n7956, CK => CLK, RN => 
                           n3072, Q => REGISTERS_51_24_port, QN => n_1547);
   REGISTERS_reg_51_23_inst : DFFR_X1 port map( D => n7957, CK => CLK, RN => 
                           n3072, Q => REGISTERS_51_23_port, QN => n_1548);
   REGISTERS_reg_51_22_inst : DFFR_X1 port map( D => n7958, CK => CLK, RN => 
                           n3072, Q => REGISTERS_51_22_port, QN => n_1549);
   REGISTERS_reg_51_21_inst : DFFR_X1 port map( D => n7959, CK => CLK, RN => 
                           n3072, Q => REGISTERS_51_21_port, QN => n_1550);
   REGISTERS_reg_51_20_inst : DFFR_X1 port map( D => n7960, CK => CLK, RN => 
                           n3072, Q => REGISTERS_51_20_port, QN => n_1551);
   REGISTERS_reg_51_19_inst : DFFR_X1 port map( D => n7961, CK => CLK, RN => 
                           n3072, Q => REGISTERS_51_19_port, QN => n_1552);
   REGISTERS_reg_51_18_inst : DFFR_X1 port map( D => n7962, CK => CLK, RN => 
                           n3072, Q => REGISTERS_51_18_port, QN => n_1553);
   REGISTERS_reg_51_17_inst : DFFR_X1 port map( D => n7963, CK => CLK, RN => 
                           n3072, Q => REGISTERS_51_17_port, QN => n_1554);
   REGISTERS_reg_51_16_inst : DFFR_X1 port map( D => n7964, CK => CLK, RN => 
                           n3072, Q => REGISTERS_51_16_port, QN => n_1555);
   REGISTERS_reg_51_15_inst : DFFR_X1 port map( D => n7965, CK => CLK, RN => 
                           n3071, Q => REGISTERS_51_15_port, QN => n_1556);
   REGISTERS_reg_51_14_inst : DFFR_X1 port map( D => n7966, CK => CLK, RN => 
                           n3071, Q => REGISTERS_51_14_port, QN => n_1557);
   REGISTERS_reg_51_13_inst : DFFR_X1 port map( D => n7967, CK => CLK, RN => 
                           n3071, Q => REGISTERS_51_13_port, QN => n_1558);
   REGISTERS_reg_51_12_inst : DFFR_X1 port map( D => n7968, CK => CLK, RN => 
                           n3071, Q => REGISTERS_51_12_port, QN => n_1559);
   REGISTERS_reg_51_11_inst : DFFR_X1 port map( D => n7969, CK => CLK, RN => 
                           n3071, Q => REGISTERS_51_11_port, QN => n_1560);
   REGISTERS_reg_51_10_inst : DFFR_X1 port map( D => n7970, CK => CLK, RN => 
                           n3071, Q => REGISTERS_51_10_port, QN => n_1561);
   REGISTERS_reg_51_9_inst : DFFR_X1 port map( D => n7971, CK => CLK, RN => 
                           n3071, Q => REGISTERS_51_9_port, QN => n_1562);
   REGISTERS_reg_51_8_inst : DFFR_X1 port map( D => n7972, CK => CLK, RN => 
                           n3071, Q => REGISTERS_51_8_port, QN => n_1563);
   REGISTERS_reg_51_7_inst : DFFR_X1 port map( D => n7973, CK => CLK, RN => 
                           n3071, Q => REGISTERS_51_7_port, QN => n_1564);
   REGISTERS_reg_51_6_inst : DFFR_X1 port map( D => n7974, CK => CLK, RN => 
                           n3071, Q => REGISTERS_51_6_port, QN => n_1565);
   REGISTERS_reg_51_5_inst : DFFR_X1 port map( D => n7975, CK => CLK, RN => 
                           n3071, Q => REGISTERS_51_5_port, QN => n_1566);
   REGISTERS_reg_51_4_inst : DFFR_X1 port map( D => n7976, CK => CLK, RN => 
                           n3071, Q => REGISTERS_51_4_port, QN => n_1567);
   REGISTERS_reg_51_3_inst : DFFR_X1 port map( D => n7977, CK => CLK, RN => 
                           n3069, Q => REGISTERS_51_3_port, QN => n_1568);
   REGISTERS_reg_51_2_inst : DFFR_X1 port map( D => n7978, CK => CLK, RN => 
                           n3069, Q => REGISTERS_51_2_port, QN => n_1569);
   REGISTERS_reg_51_1_inst : DFFR_X1 port map( D => n7979, CK => CLK, RN => 
                           n3069, Q => REGISTERS_51_1_port, QN => n_1570);
   REGISTERS_reg_51_0_inst : DFFR_X1 port map( D => n7980, CK => CLK, RN => 
                           n3069, Q => REGISTERS_51_0_port, QN => n_1571);
   REGISTERS_reg_50_31_inst : DFFR_X1 port map( D => n7917, CK => CLK, RN => 
                           n3077, Q => REGISTERS_50_31_port, QN => n_1572);
   REGISTERS_reg_50_30_inst : DFFR_X1 port map( D => n7918, CK => CLK, RN => 
                           n3077, Q => REGISTERS_50_30_port, QN => n_1573);
   REGISTERS_reg_50_29_inst : DFFR_X1 port map( D => n7919, CK => CLK, RN => 
                           n3077, Q => REGISTERS_50_29_port, QN => n_1574);
   REGISTERS_reg_50_28_inst : DFFR_X1 port map( D => n7920, CK => CLK, RN => 
                           n3077, Q => REGISTERS_50_28_port, QN => n_1575);
   REGISTERS_reg_50_27_inst : DFFR_X1 port map( D => n7921, CK => CLK, RN => 
                           n3077, Q => REGISTERS_50_27_port, QN => n_1576);
   REGISTERS_reg_50_26_inst : DFFR_X1 port map( D => n7922, CK => CLK, RN => 
                           n3077, Q => REGISTERS_50_26_port, QN => n_1577);
   REGISTERS_reg_50_25_inst : DFFR_X1 port map( D => n7923, CK => CLK, RN => 
                           n3077, Q => REGISTERS_50_25_port, QN => n_1578);
   REGISTERS_reg_50_24_inst : DFFR_X1 port map( D => n7924, CK => CLK, RN => 
                           n3077, Q => REGISTERS_50_24_port, QN => n_1579);
   REGISTERS_reg_50_23_inst : DFFR_X1 port map( D => n7925, CK => CLK, RN => 
                           n3077, Q => REGISTERS_50_23_port, QN => n_1580);
   REGISTERS_reg_50_22_inst : DFFR_X1 port map( D => n7926, CK => CLK, RN => 
                           n3077, Q => REGISTERS_50_22_port, QN => n_1581);
   REGISTERS_reg_50_21_inst : DFFR_X1 port map( D => n7927, CK => CLK, RN => 
                           n3077, Q => REGISTERS_50_21_port, QN => n_1582);
   REGISTERS_reg_50_20_inst : DFFR_X1 port map( D => n7928, CK => CLK, RN => 
                           n3077, Q => REGISTERS_50_20_port, QN => n_1583);
   REGISTERS_reg_50_19_inst : DFFR_X1 port map( D => n7929, CK => CLK, RN => 
                           n3076, Q => REGISTERS_50_19_port, QN => n_1584);
   REGISTERS_reg_50_18_inst : DFFR_X1 port map( D => n7930, CK => CLK, RN => 
                           n3076, Q => REGISTERS_50_18_port, QN => n_1585);
   REGISTERS_reg_50_17_inst : DFFR_X1 port map( D => n7931, CK => CLK, RN => 
                           n3076, Q => REGISTERS_50_17_port, QN => n_1586);
   REGISTERS_reg_50_16_inst : DFFR_X1 port map( D => n7932, CK => CLK, RN => 
                           n3076, Q => REGISTERS_50_16_port, QN => n_1587);
   REGISTERS_reg_50_15_inst : DFFR_X1 port map( D => n7933, CK => CLK, RN => 
                           n3076, Q => REGISTERS_50_15_port, QN => n_1588);
   REGISTERS_reg_50_14_inst : DFFR_X1 port map( D => n7934, CK => CLK, RN => 
                           n3076, Q => REGISTERS_50_14_port, QN => n_1589);
   REGISTERS_reg_50_13_inst : DFFR_X1 port map( D => n7935, CK => CLK, RN => 
                           n3076, Q => REGISTERS_50_13_port, QN => n_1590);
   REGISTERS_reg_50_12_inst : DFFR_X1 port map( D => n7936, CK => CLK, RN => 
                           n3076, Q => REGISTERS_50_12_port, QN => n_1591);
   REGISTERS_reg_50_11_inst : DFFR_X1 port map( D => n7937, CK => CLK, RN => 
                           n3076, Q => REGISTERS_50_11_port, QN => n_1592);
   REGISTERS_reg_50_10_inst : DFFR_X1 port map( D => n7938, CK => CLK, RN => 
                           n3076, Q => REGISTERS_50_10_port, QN => n_1593);
   REGISTERS_reg_50_9_inst : DFFR_X1 port map( D => n7939, CK => CLK, RN => 
                           n3076, Q => REGISTERS_50_9_port, QN => n_1594);
   REGISTERS_reg_50_8_inst : DFFR_X1 port map( D => n7940, CK => CLK, RN => 
                           n3076, Q => REGISTERS_50_8_port, QN => n_1595);
   REGISTERS_reg_50_7_inst : DFFR_X1 port map( D => n7941, CK => CLK, RN => 
                           n3074, Q => REGISTERS_50_7_port, QN => n_1596);
   REGISTERS_reg_50_6_inst : DFFR_X1 port map( D => n7942, CK => CLK, RN => 
                           n3074, Q => REGISTERS_50_6_port, QN => n_1597);
   REGISTERS_reg_50_5_inst : DFFR_X1 port map( D => n7943, CK => CLK, RN => 
                           n3074, Q => REGISTERS_50_5_port, QN => n_1598);
   REGISTERS_reg_50_4_inst : DFFR_X1 port map( D => n7944, CK => CLK, RN => 
                           n3074, Q => REGISTERS_50_4_port, QN => n_1599);
   REGISTERS_reg_50_3_inst : DFFR_X1 port map( D => n7945, CK => CLK, RN => 
                           n3074, Q => REGISTERS_50_3_port, QN => n_1600);
   REGISTERS_reg_50_2_inst : DFFR_X1 port map( D => n7946, CK => CLK, RN => 
                           n3074, Q => REGISTERS_50_2_port, QN => n_1601);
   REGISTERS_reg_50_1_inst : DFFR_X1 port map( D => n7947, CK => CLK, RN => 
                           n3074, Q => REGISTERS_50_1_port, QN => n_1602);
   REGISTERS_reg_50_0_inst : DFFR_X1 port map( D => n7948, CK => CLK, RN => 
                           n3074, Q => REGISTERS_50_0_port, QN => n_1603);
   REGISTERS_reg_49_31_inst : DFFR_X1 port map( D => n7885, CK => CLK, RN => 
                           n3082, Q => REGISTERS_49_31_port, QN => n_1604);
   REGISTERS_reg_49_30_inst : DFFR_X1 port map( D => n7886, CK => CLK, RN => 
                           n3082, Q => REGISTERS_49_30_port, QN => n_1605);
   REGISTERS_reg_49_29_inst : DFFR_X1 port map( D => n7887, CK => CLK, RN => 
                           n3082, Q => REGISTERS_49_29_port, QN => n_1606);
   REGISTERS_reg_49_28_inst : DFFR_X1 port map( D => n7888, CK => CLK, RN => 
                           n3082, Q => REGISTERS_49_28_port, QN => n_1607);
   REGISTERS_reg_49_27_inst : DFFR_X1 port map( D => n7889, CK => CLK, RN => 
                           n3082, Q => REGISTERS_49_27_port, QN => n_1608);
   REGISTERS_reg_49_26_inst : DFFR_X1 port map( D => n7890, CK => CLK, RN => 
                           n3082, Q => REGISTERS_49_26_port, QN => n_1609);
   REGISTERS_reg_49_25_inst : DFFR_X1 port map( D => n7891, CK => CLK, RN => 
                           n3082, Q => REGISTERS_49_25_port, QN => n_1610);
   REGISTERS_reg_49_24_inst : DFFR_X1 port map( D => n7892, CK => CLK, RN => 
                           n3082, Q => REGISTERS_49_24_port, QN => n_1611);
   REGISTERS_reg_49_23_inst : DFFR_X1 port map( D => n7893, CK => CLK, RN => 
                           n3081, Q => REGISTERS_49_23_port, QN => n_1612);
   REGISTERS_reg_49_22_inst : DFFR_X1 port map( D => n7894, CK => CLK, RN => 
                           n3081, Q => REGISTERS_49_22_port, QN => n_1613);
   REGISTERS_reg_49_21_inst : DFFR_X1 port map( D => n7895, CK => CLK, RN => 
                           n3081, Q => REGISTERS_49_21_port, QN => n_1614);
   REGISTERS_reg_49_20_inst : DFFR_X1 port map( D => n7896, CK => CLK, RN => 
                           n3081, Q => REGISTERS_49_20_port, QN => n_1615);
   REGISTERS_reg_49_19_inst : DFFR_X1 port map( D => n7897, CK => CLK, RN => 
                           n3081, Q => REGISTERS_49_19_port, QN => n_1616);
   REGISTERS_reg_49_18_inst : DFFR_X1 port map( D => n7898, CK => CLK, RN => 
                           n3081, Q => REGISTERS_49_18_port, QN => n_1617);
   REGISTERS_reg_49_17_inst : DFFR_X1 port map( D => n7899, CK => CLK, RN => 
                           n3081, Q => REGISTERS_49_17_port, QN => n_1618);
   REGISTERS_reg_49_16_inst : DFFR_X1 port map( D => n7900, CK => CLK, RN => 
                           n3081, Q => REGISTERS_49_16_port, QN => n_1619);
   REGISTERS_reg_49_15_inst : DFFR_X1 port map( D => n7901, CK => CLK, RN => 
                           n3081, Q => REGISTERS_49_15_port, QN => n_1620);
   REGISTERS_reg_49_14_inst : DFFR_X1 port map( D => n7902, CK => CLK, RN => 
                           n3081, Q => REGISTERS_49_14_port, QN => n_1621);
   REGISTERS_reg_49_13_inst : DFFR_X1 port map( D => n7903, CK => CLK, RN => 
                           n3081, Q => REGISTERS_49_13_port, QN => n_1622);
   REGISTERS_reg_49_12_inst : DFFR_X1 port map( D => n7904, CK => CLK, RN => 
                           n3081, Q => REGISTERS_49_12_port, QN => n_1623);
   REGISTERS_reg_49_11_inst : DFFR_X1 port map( D => n7905, CK => CLK, RN => 
                           n3079, Q => REGISTERS_49_11_port, QN => n_1624);
   REGISTERS_reg_49_10_inst : DFFR_X1 port map( D => n7906, CK => CLK, RN => 
                           n3079, Q => REGISTERS_49_10_port, QN => n_1625);
   REGISTERS_reg_49_9_inst : DFFR_X1 port map( D => n7907, CK => CLK, RN => 
                           n3079, Q => REGISTERS_49_9_port, QN => n_1626);
   REGISTERS_reg_49_8_inst : DFFR_X1 port map( D => n7908, CK => CLK, RN => 
                           n3079, Q => REGISTERS_49_8_port, QN => n_1627);
   REGISTERS_reg_49_7_inst : DFFR_X1 port map( D => n7909, CK => CLK, RN => 
                           n3079, Q => REGISTERS_49_7_port, QN => n_1628);
   REGISTERS_reg_49_6_inst : DFFR_X1 port map( D => n7910, CK => CLK, RN => 
                           n3079, Q => REGISTERS_49_6_port, QN => n_1629);
   REGISTERS_reg_49_5_inst : DFFR_X1 port map( D => n7911, CK => CLK, RN => 
                           n3079, Q => REGISTERS_49_5_port, QN => n_1630);
   REGISTERS_reg_49_4_inst : DFFR_X1 port map( D => n7912, CK => CLK, RN => 
                           n3079, Q => REGISTERS_49_4_port, QN => n_1631);
   REGISTERS_reg_49_3_inst : DFFR_X1 port map( D => n7913, CK => CLK, RN => 
                           n3079, Q => REGISTERS_49_3_port, QN => n_1632);
   REGISTERS_reg_49_2_inst : DFFR_X1 port map( D => n7914, CK => CLK, RN => 
                           n3079, Q => REGISTERS_49_2_port, QN => n_1633);
   REGISTERS_reg_49_1_inst : DFFR_X1 port map( D => n7915, CK => CLK, RN => 
                           n3079, Q => REGISTERS_49_1_port, QN => n_1634);
   REGISTERS_reg_49_0_inst : DFFR_X1 port map( D => n7916, CK => CLK, RN => 
                           n3079, Q => REGISTERS_49_0_port, QN => n_1635);
   REGISTERS_reg_45_31_inst : DFFR_X1 port map( D => n7757, CK => CLK, RN => 
                           n3101, Q => REGISTERS_45_31_port, QN => n_1636);
   REGISTERS_reg_45_30_inst : DFFR_X1 port map( D => n7758, CK => CLK, RN => 
                           n3101, Q => REGISTERS_45_30_port, QN => n_1637);
   REGISTERS_reg_45_29_inst : DFFR_X1 port map( D => n7759, CK => CLK, RN => 
                           n3101, Q => REGISTERS_45_29_port, QN => n_1638);
   REGISTERS_reg_45_28_inst : DFFR_X1 port map( D => n7760, CK => CLK, RN => 
                           n3101, Q => REGISTERS_45_28_port, QN => n_1639);
   REGISTERS_reg_45_27_inst : DFFR_X1 port map( D => n7761, CK => CLK, RN => 
                           n3099, Q => REGISTERS_45_27_port, QN => n_1640);
   REGISTERS_reg_45_26_inst : DFFR_X1 port map( D => n7762, CK => CLK, RN => 
                           n3099, Q => REGISTERS_45_26_port, QN => n_1641);
   REGISTERS_reg_45_25_inst : DFFR_X1 port map( D => n7763, CK => CLK, RN => 
                           n3099, Q => REGISTERS_45_25_port, QN => n_1642);
   REGISTERS_reg_45_24_inst : DFFR_X1 port map( D => n7764, CK => CLK, RN => 
                           n3099, Q => REGISTERS_45_24_port, QN => n_1643);
   REGISTERS_reg_45_23_inst : DFFR_X1 port map( D => n7765, CK => CLK, RN => 
                           n3099, Q => REGISTERS_45_23_port, QN => n_1644);
   REGISTERS_reg_45_22_inst : DFFR_X1 port map( D => n7766, CK => CLK, RN => 
                           n3099, Q => REGISTERS_45_22_port, QN => n_1645);
   REGISTERS_reg_45_21_inst : DFFR_X1 port map( D => n7767, CK => CLK, RN => 
                           n3099, Q => REGISTERS_45_21_port, QN => n_1646);
   REGISTERS_reg_45_20_inst : DFFR_X1 port map( D => n7768, CK => CLK, RN => 
                           n3099, Q => REGISTERS_45_20_port, QN => n_1647);
   REGISTERS_reg_45_19_inst : DFFR_X1 port map( D => n7769, CK => CLK, RN => 
                           n3099, Q => REGISTERS_45_19_port, QN => n_1648);
   REGISTERS_reg_45_18_inst : DFFR_X1 port map( D => n7770, CK => CLK, RN => 
                           n3099, Q => REGISTERS_45_18_port, QN => n_1649);
   REGISTERS_reg_45_17_inst : DFFR_X1 port map( D => n7771, CK => CLK, RN => 
                           n3099, Q => REGISTERS_45_17_port, QN => n_1650);
   REGISTERS_reg_45_16_inst : DFFR_X1 port map( D => n7772, CK => CLK, RN => 
                           n3099, Q => REGISTERS_45_16_port, QN => n_1651);
   REGISTERS_reg_45_15_inst : DFFR_X1 port map( D => n7773, CK => CLK, RN => 
                           n3097, Q => REGISTERS_45_15_port, QN => n_1652);
   REGISTERS_reg_45_14_inst : DFFR_X1 port map( D => n7774, CK => CLK, RN => 
                           n3097, Q => REGISTERS_45_14_port, QN => n_1653);
   REGISTERS_reg_45_13_inst : DFFR_X1 port map( D => n7775, CK => CLK, RN => 
                           n3097, Q => REGISTERS_45_13_port, QN => n_1654);
   REGISTERS_reg_45_12_inst : DFFR_X1 port map( D => n7776, CK => CLK, RN => 
                           n3097, Q => REGISTERS_45_12_port, QN => n_1655);
   REGISTERS_reg_45_11_inst : DFFR_X1 port map( D => n7777, CK => CLK, RN => 
                           n3097, Q => REGISTERS_45_11_port, QN => n_1656);
   REGISTERS_reg_45_10_inst : DFFR_X1 port map( D => n7778, CK => CLK, RN => 
                           n3097, Q => REGISTERS_45_10_port, QN => n_1657);
   REGISTERS_reg_45_9_inst : DFFR_X1 port map( D => n7779, CK => CLK, RN => 
                           n3097, Q => REGISTERS_45_9_port, QN => n_1658);
   REGISTERS_reg_45_8_inst : DFFR_X1 port map( D => n7780, CK => CLK, RN => 
                           n3097, Q => REGISTERS_45_8_port, QN => n_1659);
   REGISTERS_reg_45_7_inst : DFFR_X1 port map( D => n7781, CK => CLK, RN => 
                           n3097, Q => REGISTERS_45_7_port, QN => n_1660);
   REGISTERS_reg_45_6_inst : DFFR_X1 port map( D => n7782, CK => CLK, RN => 
                           n3097, Q => REGISTERS_45_6_port, QN => n_1661);
   REGISTERS_reg_45_5_inst : DFFR_X1 port map( D => n7783, CK => CLK, RN => 
                           n3097, Q => REGISTERS_45_5_port, QN => n_1662);
   REGISTERS_reg_45_4_inst : DFFR_X1 port map( D => n7784, CK => CLK, RN => 
                           n3097, Q => REGISTERS_45_4_port, QN => n_1663);
   REGISTERS_reg_45_3_inst : DFFR_X1 port map( D => n7785, CK => CLK, RN => 
                           n3096, Q => REGISTERS_45_3_port, QN => n_1664);
   REGISTERS_reg_45_2_inst : DFFR_X1 port map( D => n7786, CK => CLK, RN => 
                           n3096, Q => REGISTERS_45_2_port, QN => n_1665);
   REGISTERS_reg_45_1_inst : DFFR_X1 port map( D => n7787, CK => CLK, RN => 
                           n3096, Q => REGISTERS_45_1_port, QN => n_1666);
   REGISTERS_reg_45_0_inst : DFFR_X1 port map( D => n7788, CK => CLK, RN => 
                           n3096, Q => REGISTERS_45_0_port, QN => n_1667);
   REGISTERS_reg_44_31_inst : DFFR_X1 port map( D => n7725, CK => CLK, RN => 
                           n3104, Q => REGISTERS_44_31_port, QN => n_1668);
   REGISTERS_reg_44_30_inst : DFFR_X1 port map( D => n7726, CK => CLK, RN => 
                           n3104, Q => REGISTERS_44_30_port, QN => n_1669);
   REGISTERS_reg_44_29_inst : DFFR_X1 port map( D => n7727, CK => CLK, RN => 
                           n3104, Q => REGISTERS_44_29_port, QN => n_1670);
   REGISTERS_reg_44_28_inst : DFFR_X1 port map( D => n7728, CK => CLK, RN => 
                           n3104, Q => REGISTERS_44_28_port, QN => n_1671);
   REGISTERS_reg_44_27_inst : DFFR_X1 port map( D => n7729, CK => CLK, RN => 
                           n3104, Q => REGISTERS_44_27_port, QN => n_1672);
   REGISTERS_reg_44_26_inst : DFFR_X1 port map( D => n7730, CK => CLK, RN => 
                           n3104, Q => REGISTERS_44_26_port, QN => n_1673);
   REGISTERS_reg_44_25_inst : DFFR_X1 port map( D => n7731, CK => CLK, RN => 
                           n3104, Q => REGISTERS_44_25_port, QN => n_1674);
   REGISTERS_reg_44_24_inst : DFFR_X1 port map( D => n7732, CK => CLK, RN => 
                           n3104, Q => REGISTERS_44_24_port, QN => n_1675);
   REGISTERS_reg_44_23_inst : DFFR_X1 port map( D => n7733, CK => CLK, RN => 
                           n3104, Q => REGISTERS_44_23_port, QN => n_1676);
   REGISTERS_reg_44_22_inst : DFFR_X1 port map( D => n7734, CK => CLK, RN => 
                           n3104, Q => REGISTERS_44_22_port, QN => n_1677);
   REGISTERS_reg_44_21_inst : DFFR_X1 port map( D => n7735, CK => CLK, RN => 
                           n3104, Q => REGISTERS_44_21_port, QN => n_1678);
   REGISTERS_reg_44_20_inst : DFFR_X1 port map( D => n7736, CK => CLK, RN => 
                           n3104, Q => REGISTERS_44_20_port, QN => n_1679);
   REGISTERS_reg_44_19_inst : DFFR_X1 port map( D => n7737, CK => CLK, RN => 
                           n3102, Q => REGISTERS_44_19_port, QN => n_1680);
   REGISTERS_reg_44_18_inst : DFFR_X1 port map( D => n7738, CK => CLK, RN => 
                           n3102, Q => REGISTERS_44_18_port, QN => n_1681);
   REGISTERS_reg_44_17_inst : DFFR_X1 port map( D => n7739, CK => CLK, RN => 
                           n3102, Q => REGISTERS_44_17_port, QN => n_1682);
   REGISTERS_reg_44_16_inst : DFFR_X1 port map( D => n7740, CK => CLK, RN => 
                           n3102, Q => REGISTERS_44_16_port, QN => n_1683);
   REGISTERS_reg_44_15_inst : DFFR_X1 port map( D => n7741, CK => CLK, RN => 
                           n3102, Q => REGISTERS_44_15_port, QN => n_1684);
   REGISTERS_reg_44_14_inst : DFFR_X1 port map( D => n7742, CK => CLK, RN => 
                           n3102, Q => REGISTERS_44_14_port, QN => n_1685);
   REGISTERS_reg_44_13_inst : DFFR_X1 port map( D => n7743, CK => CLK, RN => 
                           n3102, Q => REGISTERS_44_13_port, QN => n_1686);
   REGISTERS_reg_44_12_inst : DFFR_X1 port map( D => n7744, CK => CLK, RN => 
                           n3102, Q => REGISTERS_44_12_port, QN => n_1687);
   REGISTERS_reg_44_11_inst : DFFR_X1 port map( D => n7745, CK => CLK, RN => 
                           n3102, Q => REGISTERS_44_11_port, QN => n_1688);
   REGISTERS_reg_44_10_inst : DFFR_X1 port map( D => n7746, CK => CLK, RN => 
                           n3102, Q => REGISTERS_44_10_port, QN => n_1689);
   REGISTERS_reg_44_9_inst : DFFR_X1 port map( D => n7747, CK => CLK, RN => 
                           n3102, Q => REGISTERS_44_9_port, QN => n_1690);
   REGISTERS_reg_44_8_inst : DFFR_X1 port map( D => n7748, CK => CLK, RN => 
                           n3102, Q => REGISTERS_44_8_port, QN => n_1691);
   REGISTERS_reg_44_7_inst : DFFR_X1 port map( D => n7749, CK => CLK, RN => 
                           n3101, Q => REGISTERS_44_7_port, QN => n_1692);
   REGISTERS_reg_44_6_inst : DFFR_X1 port map( D => n7750, CK => CLK, RN => 
                           n3101, Q => REGISTERS_44_6_port, QN => n_1693);
   REGISTERS_reg_44_5_inst : DFFR_X1 port map( D => n7751, CK => CLK, RN => 
                           n3101, Q => REGISTERS_44_5_port, QN => n_1694);
   REGISTERS_reg_44_4_inst : DFFR_X1 port map( D => n7752, CK => CLK, RN => 
                           n3101, Q => REGISTERS_44_4_port, QN => n_1695);
   REGISTERS_reg_44_3_inst : DFFR_X1 port map( D => n7753, CK => CLK, RN => 
                           n3101, Q => REGISTERS_44_3_port, QN => n_1696);
   REGISTERS_reg_44_2_inst : DFFR_X1 port map( D => n7754, CK => CLK, RN => 
                           n3101, Q => REGISTERS_44_2_port, QN => n_1697);
   REGISTERS_reg_44_1_inst : DFFR_X1 port map( D => n7755, CK => CLK, RN => 
                           n3101, Q => REGISTERS_44_1_port, QN => n_1698);
   REGISTERS_reg_44_0_inst : DFFR_X1 port map( D => n7756, CK => CLK, RN => 
                           n3101, Q => REGISTERS_44_0_port, QN => n_1699);
   REGISTERS_reg_43_31_inst : DFFR_X1 port map( D => n7693, CK => CLK, RN => 
                           n3113, Q => REGISTERS_43_31_port, QN => n_1700);
   REGISTERS_reg_43_30_inst : DFFR_X1 port map( D => n7694, CK => CLK, RN => 
                           n3113, Q => REGISTERS_43_30_port, QN => n_1701);
   REGISTERS_reg_43_29_inst : DFFR_X1 port map( D => n7695, CK => CLK, RN => 
                           n3113, Q => REGISTERS_43_29_port, QN => n_1702);
   REGISTERS_reg_43_28_inst : DFFR_X1 port map( D => n7696, CK => CLK, RN => 
                           n3113, Q => REGISTERS_43_28_port, QN => n_1703);
   REGISTERS_reg_43_27_inst : DFFR_X1 port map( D => n7697, CK => CLK, RN => 
                           n3113, Q => REGISTERS_43_27_port, QN => n_1704);
   REGISTERS_reg_43_26_inst : DFFR_X1 port map( D => n7698, CK => CLK, RN => 
                           n3113, Q => REGISTERS_43_26_port, QN => n_1705);
   REGISTERS_reg_43_25_inst : DFFR_X1 port map( D => n7699, CK => CLK, RN => 
                           n3113, Q => REGISTERS_43_25_port, QN => n_1706);
   REGISTERS_reg_43_24_inst : DFFR_X1 port map( D => n7700, CK => CLK, RN => 
                           n3113, Q => REGISTERS_43_24_port, QN => n_1707);
   REGISTERS_reg_43_23_inst : DFFR_X1 port map( D => n7701, CK => CLK, RN => 
                           n3111, Q => REGISTERS_43_23_port, QN => n_1708);
   REGISTERS_reg_43_22_inst : DFFR_X1 port map( D => n7702, CK => CLK, RN => 
                           n3111, Q => REGISTERS_43_22_port, QN => n_1709);
   REGISTERS_reg_43_21_inst : DFFR_X1 port map( D => n7703, CK => CLK, RN => 
                           n3111, Q => REGISTERS_43_21_port, QN => n_1710);
   REGISTERS_reg_43_20_inst : DFFR_X1 port map( D => n7704, CK => CLK, RN => 
                           n3111, Q => REGISTERS_43_20_port, QN => n_1711);
   REGISTERS_reg_43_19_inst : DFFR_X1 port map( D => n7705, CK => CLK, RN => 
                           n3111, Q => REGISTERS_43_19_port, QN => n_1712);
   REGISTERS_reg_43_18_inst : DFFR_X1 port map( D => n7706, CK => CLK, RN => 
                           n3111, Q => REGISTERS_43_18_port, QN => n_1713);
   REGISTERS_reg_43_17_inst : DFFR_X1 port map( D => n7707, CK => CLK, RN => 
                           n3111, Q => REGISTERS_43_17_port, QN => n_1714);
   REGISTERS_reg_43_16_inst : DFFR_X1 port map( D => n7708, CK => CLK, RN => 
                           n3111, Q => REGISTERS_43_16_port, QN => n_1715);
   REGISTERS_reg_43_15_inst : DFFR_X1 port map( D => n7709, CK => CLK, RN => 
                           n3111, Q => REGISTERS_43_15_port, QN => n_1716);
   REGISTERS_reg_43_14_inst : DFFR_X1 port map( D => n7710, CK => CLK, RN => 
                           n3111, Q => REGISTERS_43_14_port, QN => n_1717);
   REGISTERS_reg_43_13_inst : DFFR_X1 port map( D => n7711, CK => CLK, RN => 
                           n3111, Q => REGISTERS_43_13_port, QN => n_1718);
   REGISTERS_reg_43_12_inst : DFFR_X1 port map( D => n7712, CK => CLK, RN => 
                           n3111, Q => REGISTERS_43_12_port, QN => n_1719);
   REGISTERS_reg_43_11_inst : DFFR_X1 port map( D => n7713, CK => CLK, RN => 
                           n3110, Q => REGISTERS_43_11_port, QN => n_1720);
   REGISTERS_reg_43_10_inst : DFFR_X1 port map( D => n7714, CK => CLK, RN => 
                           n3110, Q => REGISTERS_43_10_port, QN => n_1721);
   REGISTERS_reg_43_9_inst : DFFR_X1 port map( D => n7715, CK => CLK, RN => 
                           n3110, Q => REGISTERS_43_9_port, QN => n_1722);
   REGISTERS_reg_43_8_inst : DFFR_X1 port map( D => n7716, CK => CLK, RN => 
                           n3110, Q => REGISTERS_43_8_port, QN => n_1723);
   REGISTERS_reg_43_7_inst : DFFR_X1 port map( D => n7717, CK => CLK, RN => 
                           n3110, Q => REGISTERS_43_7_port, QN => n_1724);
   REGISTERS_reg_43_6_inst : DFFR_X1 port map( D => n7718, CK => CLK, RN => 
                           n3110, Q => REGISTERS_43_6_port, QN => n_1725);
   REGISTERS_reg_43_5_inst : DFFR_X1 port map( D => n7719, CK => CLK, RN => 
                           n3110, Q => REGISTERS_43_5_port, QN => n_1726);
   REGISTERS_reg_43_4_inst : DFFR_X1 port map( D => n7720, CK => CLK, RN => 
                           n3110, Q => REGISTERS_43_4_port, QN => n_1727);
   REGISTERS_reg_43_3_inst : DFFR_X1 port map( D => n7721, CK => CLK, RN => 
                           n3110, Q => REGISTERS_43_3_port, QN => n_1728);
   REGISTERS_reg_43_2_inst : DFFR_X1 port map( D => n7722, CK => CLK, RN => 
                           n3110, Q => REGISTERS_43_2_port, QN => n_1729);
   REGISTERS_reg_43_1_inst : DFFR_X1 port map( D => n7723, CK => CLK, RN => 
                           n3110, Q => REGISTERS_43_1_port, QN => n_1730);
   REGISTERS_reg_43_0_inst : DFFR_X1 port map( D => n7724, CK => CLK, RN => 
                           n3110, Q => REGISTERS_43_0_port, QN => n_1731);
   REGISTERS_reg_42_31_inst : DFFR_X1 port map( D => n7661, CK => CLK, RN => 
                           n3118, Q => REGISTERS_42_31_port, QN => n_1732);
   REGISTERS_reg_42_30_inst : DFFR_X1 port map( D => n7662, CK => CLK, RN => 
                           n3118, Q => REGISTERS_42_30_port, QN => n_1733);
   REGISTERS_reg_42_29_inst : DFFR_X1 port map( D => n7663, CK => CLK, RN => 
                           n3118, Q => REGISTERS_42_29_port, QN => n_1734);
   REGISTERS_reg_42_28_inst : DFFR_X1 port map( D => n7664, CK => CLK, RN => 
                           n3118, Q => REGISTERS_42_28_port, QN => n_1735);
   REGISTERS_reg_42_27_inst : DFFR_X1 port map( D => n7665, CK => CLK, RN => 
                           n3116, Q => REGISTERS_42_27_port, QN => n_1736);
   REGISTERS_reg_42_26_inst : DFFR_X1 port map( D => n7666, CK => CLK, RN => 
                           n3116, Q => REGISTERS_42_26_port, QN => n_1737);
   REGISTERS_reg_42_25_inst : DFFR_X1 port map( D => n7667, CK => CLK, RN => 
                           n3116, Q => REGISTERS_42_25_port, QN => n_1738);
   REGISTERS_reg_42_24_inst : DFFR_X1 port map( D => n7668, CK => CLK, RN => 
                           n3116, Q => REGISTERS_42_24_port, QN => n_1739);
   REGISTERS_reg_42_23_inst : DFFR_X1 port map( D => n7669, CK => CLK, RN => 
                           n3116, Q => REGISTERS_42_23_port, QN => n_1740);
   REGISTERS_reg_42_22_inst : DFFR_X1 port map( D => n7670, CK => CLK, RN => 
                           n3116, Q => REGISTERS_42_22_port, QN => n_1741);
   REGISTERS_reg_42_21_inst : DFFR_X1 port map( D => n7671, CK => CLK, RN => 
                           n3116, Q => REGISTERS_42_21_port, QN => n_1742);
   REGISTERS_reg_42_20_inst : DFFR_X1 port map( D => n7672, CK => CLK, RN => 
                           n3116, Q => REGISTERS_42_20_port, QN => n_1743);
   REGISTERS_reg_42_19_inst : DFFR_X1 port map( D => n7673, CK => CLK, RN => 
                           n3116, Q => REGISTERS_42_19_port, QN => n_1744);
   REGISTERS_reg_42_18_inst : DFFR_X1 port map( D => n7674, CK => CLK, RN => 
                           n3116, Q => REGISTERS_42_18_port, QN => n_1745);
   REGISTERS_reg_42_17_inst : DFFR_X1 port map( D => n7675, CK => CLK, RN => 
                           n3116, Q => REGISTERS_42_17_port, QN => n_1746);
   REGISTERS_reg_42_16_inst : DFFR_X1 port map( D => n7676, CK => CLK, RN => 
                           n3116, Q => REGISTERS_42_16_port, QN => n_1747);
   REGISTERS_reg_42_15_inst : DFFR_X1 port map( D => n7677, CK => CLK, RN => 
                           n3115, Q => REGISTERS_42_15_port, QN => n_1748);
   REGISTERS_reg_42_14_inst : DFFR_X1 port map( D => n7678, CK => CLK, RN => 
                           n3115, Q => REGISTERS_42_14_port, QN => n_1749);
   REGISTERS_reg_42_13_inst : DFFR_X1 port map( D => n7679, CK => CLK, RN => 
                           n3115, Q => REGISTERS_42_13_port, QN => n_1750);
   REGISTERS_reg_42_12_inst : DFFR_X1 port map( D => n7680, CK => CLK, RN => 
                           n3115, Q => REGISTERS_42_12_port, QN => n_1751);
   REGISTERS_reg_42_11_inst : DFFR_X1 port map( D => n7681, CK => CLK, RN => 
                           n3115, Q => REGISTERS_42_11_port, QN => n_1752);
   REGISTERS_reg_42_10_inst : DFFR_X1 port map( D => n7682, CK => CLK, RN => 
                           n3115, Q => REGISTERS_42_10_port, QN => n_1753);
   REGISTERS_reg_42_9_inst : DFFR_X1 port map( D => n7683, CK => CLK, RN => 
                           n3115, Q => REGISTERS_42_9_port, QN => n_1754);
   REGISTERS_reg_42_8_inst : DFFR_X1 port map( D => n7684, CK => CLK, RN => 
                           n3115, Q => REGISTERS_42_8_port, QN => n_1755);
   REGISTERS_reg_42_7_inst : DFFR_X1 port map( D => n7685, CK => CLK, RN => 
                           n3115, Q => REGISTERS_42_7_port, QN => n_1756);
   REGISTERS_reg_42_6_inst : DFFR_X1 port map( D => n7686, CK => CLK, RN => 
                           n3115, Q => REGISTERS_42_6_port, QN => n_1757);
   REGISTERS_reg_42_5_inst : DFFR_X1 port map( D => n7687, CK => CLK, RN => 
                           n3115, Q => REGISTERS_42_5_port, QN => n_1758);
   REGISTERS_reg_42_4_inst : DFFR_X1 port map( D => n7688, CK => CLK, RN => 
                           n3115, Q => REGISTERS_42_4_port, QN => n_1759);
   REGISTERS_reg_42_3_inst : DFFR_X1 port map( D => n7689, CK => CLK, RN => 
                           n3113, Q => REGISTERS_42_3_port, QN => n_1760);
   REGISTERS_reg_42_2_inst : DFFR_X1 port map( D => n7690, CK => CLK, RN => 
                           n3113, Q => REGISTERS_42_2_port, QN => n_1761);
   REGISTERS_reg_42_1_inst : DFFR_X1 port map( D => n7691, CK => CLK, RN => 
                           n3113, Q => REGISTERS_42_1_port, QN => n_1762);
   REGISTERS_reg_42_0_inst : DFFR_X1 port map( D => n7692, CK => CLK, RN => 
                           n3113, Q => REGISTERS_42_0_port, QN => n_1763);
   REGISTERS_reg_41_31_inst : DFFR_X1 port map( D => n7629, CK => CLK, RN => 
                           n3120, Q => REGISTERS_41_31_port, QN => n_1764);
   REGISTERS_reg_41_30_inst : DFFR_X1 port map( D => n7630, CK => CLK, RN => 
                           n3120, Q => REGISTERS_41_30_port, QN => n_1765);
   REGISTERS_reg_41_29_inst : DFFR_X1 port map( D => n7631, CK => CLK, RN => 
                           n3120, Q => REGISTERS_41_29_port, QN => n_1766);
   REGISTERS_reg_41_28_inst : DFFR_X1 port map( D => n7632, CK => CLK, RN => 
                           n3120, Q => REGISTERS_41_28_port, QN => n_1767);
   REGISTERS_reg_41_27_inst : DFFR_X1 port map( D => n7633, CK => CLK, RN => 
                           n3120, Q => REGISTERS_41_27_port, QN => n_1768);
   REGISTERS_reg_41_26_inst : DFFR_X1 port map( D => n7634, CK => CLK, RN => 
                           n3120, Q => REGISTERS_41_26_port, QN => n_1769);
   REGISTERS_reg_41_25_inst : DFFR_X1 port map( D => n7635, CK => CLK, RN => 
                           n3120, Q => REGISTERS_41_25_port, QN => n_1770);
   REGISTERS_reg_41_24_inst : DFFR_X1 port map( D => n7636, CK => CLK, RN => 
                           n3120, Q => REGISTERS_41_24_port, QN => n_1771);
   REGISTERS_reg_41_23_inst : DFFR_X1 port map( D => n7637, CK => CLK, RN => 
                           n3120, Q => REGISTERS_41_23_port, QN => n_1772);
   REGISTERS_reg_41_22_inst : DFFR_X1 port map( D => n7638, CK => CLK, RN => 
                           n3120, Q => REGISTERS_41_22_port, QN => n_1773);
   REGISTERS_reg_41_21_inst : DFFR_X1 port map( D => n7639, CK => CLK, RN => 
                           n3120, Q => REGISTERS_41_21_port, QN => n_1774);
   REGISTERS_reg_41_20_inst : DFFR_X1 port map( D => n7640, CK => CLK, RN => 
                           n3120, Q => REGISTERS_41_20_port, QN => n_1775);
   REGISTERS_reg_41_19_inst : DFFR_X1 port map( D => n7641, CK => CLK, RN => 
                           n3119, Q => REGISTERS_41_19_port, QN => n_1776);
   REGISTERS_reg_41_18_inst : DFFR_X1 port map( D => n7642, CK => CLK, RN => 
                           n3119, Q => REGISTERS_41_18_port, QN => n_1777);
   REGISTERS_reg_41_17_inst : DFFR_X1 port map( D => n7643, CK => CLK, RN => 
                           n3119, Q => REGISTERS_41_17_port, QN => n_1778);
   REGISTERS_reg_41_16_inst : DFFR_X1 port map( D => n7644, CK => CLK, RN => 
                           n3119, Q => REGISTERS_41_16_port, QN => n_1779);
   REGISTERS_reg_41_15_inst : DFFR_X1 port map( D => n7645, CK => CLK, RN => 
                           n3119, Q => REGISTERS_41_15_port, QN => n_1780);
   REGISTERS_reg_41_14_inst : DFFR_X1 port map( D => n7646, CK => CLK, RN => 
                           n3119, Q => REGISTERS_41_14_port, QN => n_1781);
   REGISTERS_reg_41_13_inst : DFFR_X1 port map( D => n7647, CK => CLK, RN => 
                           n3119, Q => REGISTERS_41_13_port, QN => n_1782);
   REGISTERS_reg_41_12_inst : DFFR_X1 port map( D => n7648, CK => CLK, RN => 
                           n3119, Q => REGISTERS_41_12_port, QN => n_1783);
   REGISTERS_reg_41_11_inst : DFFR_X1 port map( D => n7649, CK => CLK, RN => 
                           n3119, Q => REGISTERS_41_11_port, QN => n_1784);
   REGISTERS_reg_41_10_inst : DFFR_X1 port map( D => n7650, CK => CLK, RN => 
                           n3119, Q => REGISTERS_41_10_port, QN => n_1785);
   REGISTERS_reg_41_9_inst : DFFR_X1 port map( D => n7651, CK => CLK, RN => 
                           n3119, Q => REGISTERS_41_9_port, QN => n_1786);
   REGISTERS_reg_41_8_inst : DFFR_X1 port map( D => n7652, CK => CLK, RN => 
                           n3119, Q => REGISTERS_41_8_port, QN => n_1787);
   REGISTERS_reg_41_7_inst : DFFR_X1 port map( D => n7653, CK => CLK, RN => 
                           n3118, Q => REGISTERS_41_7_port, QN => n_1788);
   REGISTERS_reg_41_6_inst : DFFR_X1 port map( D => n7654, CK => CLK, RN => 
                           n3118, Q => REGISTERS_41_6_port, QN => n_1789);
   REGISTERS_reg_41_5_inst : DFFR_X1 port map( D => n7655, CK => CLK, RN => 
                           n3118, Q => REGISTERS_41_5_port, QN => n_1790);
   REGISTERS_reg_41_4_inst : DFFR_X1 port map( D => n7656, CK => CLK, RN => 
                           n3118, Q => REGISTERS_41_4_port, QN => n_1791);
   REGISTERS_reg_41_3_inst : DFFR_X1 port map( D => n7657, CK => CLK, RN => 
                           n3118, Q => REGISTERS_41_3_port, QN => n_1792);
   REGISTERS_reg_41_2_inst : DFFR_X1 port map( D => n7658, CK => CLK, RN => 
                           n3118, Q => REGISTERS_41_2_port, QN => n_1793);
   REGISTERS_reg_41_1_inst : DFFR_X1 port map( D => n7659, CK => CLK, RN => 
                           n3118, Q => REGISTERS_41_1_port, QN => n_1794);
   REGISTERS_reg_41_0_inst : DFFR_X1 port map( D => n7660, CK => CLK, RN => 
                           n3118, Q => REGISTERS_41_0_port, QN => n_1795);
   REGISTERS_reg_40_31_inst : DFFR_X1 port map( D => n7597, CK => CLK, RN => 
                           n3124, Q => REGISTERS_40_31_port, QN => n_1796);
   REGISTERS_reg_40_30_inst : DFFR_X1 port map( D => n7598, CK => CLK, RN => 
                           n3124, Q => REGISTERS_40_30_port, QN => n_1797);
   REGISTERS_reg_40_29_inst : DFFR_X1 port map( D => n7599, CK => CLK, RN => 
                           n3124, Q => REGISTERS_40_29_port, QN => n_1798);
   REGISTERS_reg_40_28_inst : DFFR_X1 port map( D => n7600, CK => CLK, RN => 
                           n3124, Q => REGISTERS_40_28_port, QN => n_1799);
   REGISTERS_reg_40_27_inst : DFFR_X1 port map( D => n7601, CK => CLK, RN => 
                           n3124, Q => REGISTERS_40_27_port, QN => n_1800);
   REGISTERS_reg_40_26_inst : DFFR_X1 port map( D => n7602, CK => CLK, RN => 
                           n3124, Q => REGISTERS_40_26_port, QN => n_1801);
   REGISTERS_reg_40_25_inst : DFFR_X1 port map( D => n7603, CK => CLK, RN => 
                           n3124, Q => REGISTERS_40_25_port, QN => n_1802);
   REGISTERS_reg_40_24_inst : DFFR_X1 port map( D => n7604, CK => CLK, RN => 
                           n3124, Q => REGISTERS_40_24_port, QN => n_1803);
   REGISTERS_reg_40_23_inst : DFFR_X1 port map( D => n7605, CK => CLK, RN => 
                           n3123, Q => REGISTERS_40_23_port, QN => n_1804);
   REGISTERS_reg_40_22_inst : DFFR_X1 port map( D => n7606, CK => CLK, RN => 
                           n3123, Q => REGISTERS_40_22_port, QN => n_1805);
   REGISTERS_reg_40_21_inst : DFFR_X1 port map( D => n7607, CK => CLK, RN => 
                           n3123, Q => REGISTERS_40_21_port, QN => n_1806);
   REGISTERS_reg_40_20_inst : DFFR_X1 port map( D => n7608, CK => CLK, RN => 
                           n3123, Q => REGISTERS_40_20_port, QN => n_1807);
   REGISTERS_reg_40_19_inst : DFFR_X1 port map( D => n7609, CK => CLK, RN => 
                           n3123, Q => REGISTERS_40_19_port, QN => n_1808);
   REGISTERS_reg_40_18_inst : DFFR_X1 port map( D => n7610, CK => CLK, RN => 
                           n3123, Q => REGISTERS_40_18_port, QN => n_1809);
   REGISTERS_reg_40_17_inst : DFFR_X1 port map( D => n7611, CK => CLK, RN => 
                           n3123, Q => REGISTERS_40_17_port, QN => n_1810);
   REGISTERS_reg_40_16_inst : DFFR_X1 port map( D => n7612, CK => CLK, RN => 
                           n3123, Q => REGISTERS_40_16_port, QN => n_1811);
   REGISTERS_reg_40_15_inst : DFFR_X1 port map( D => n7613, CK => CLK, RN => 
                           n3123, Q => REGISTERS_40_15_port, QN => n_1812);
   REGISTERS_reg_40_14_inst : DFFR_X1 port map( D => n7614, CK => CLK, RN => 
                           n3123, Q => REGISTERS_40_14_port, QN => n_1813);
   REGISTERS_reg_40_13_inst : DFFR_X1 port map( D => n7615, CK => CLK, RN => 
                           n3123, Q => REGISTERS_40_13_port, QN => n_1814);
   REGISTERS_reg_40_12_inst : DFFR_X1 port map( D => n7616, CK => CLK, RN => 
                           n3123, Q => REGISTERS_40_12_port, QN => n_1815);
   REGISTERS_reg_40_11_inst : DFFR_X1 port map( D => n7617, CK => CLK, RN => 
                           n3122, Q => REGISTERS_40_11_port, QN => n_1816);
   REGISTERS_reg_40_10_inst : DFFR_X1 port map( D => n7618, CK => CLK, RN => 
                           n3122, Q => REGISTERS_40_10_port, QN => n_1817);
   REGISTERS_reg_40_9_inst : DFFR_X1 port map( D => n7619, CK => CLK, RN => 
                           n3122, Q => REGISTERS_40_9_port, QN => n_1818);
   REGISTERS_reg_40_8_inst : DFFR_X1 port map( D => n7620, CK => CLK, RN => 
                           n3122, Q => REGISTERS_40_8_port, QN => n_1819);
   REGISTERS_reg_40_7_inst : DFFR_X1 port map( D => n7621, CK => CLK, RN => 
                           n3122, Q => REGISTERS_40_7_port, QN => n_1820);
   REGISTERS_reg_40_6_inst : DFFR_X1 port map( D => n7622, CK => CLK, RN => 
                           n3122, Q => REGISTERS_40_6_port, QN => n_1821);
   REGISTERS_reg_40_5_inst : DFFR_X1 port map( D => n7623, CK => CLK, RN => 
                           n3122, Q => REGISTERS_40_5_port, QN => n_1822);
   REGISTERS_reg_40_4_inst : DFFR_X1 port map( D => n7624, CK => CLK, RN => 
                           n3122, Q => REGISTERS_40_4_port, QN => n_1823);
   REGISTERS_reg_40_3_inst : DFFR_X1 port map( D => n7625, CK => CLK, RN => 
                           n3122, Q => REGISTERS_40_3_port, QN => n_1824);
   REGISTERS_reg_40_2_inst : DFFR_X1 port map( D => n7626, CK => CLK, RN => 
                           n3122, Q => REGISTERS_40_2_port, QN => n_1825);
   REGISTERS_reg_40_1_inst : DFFR_X1 port map( D => n7627, CK => CLK, RN => 
                           n3122, Q => REGISTERS_40_1_port, QN => n_1826);
   REGISTERS_reg_40_0_inst : DFFR_X1 port map( D => n7628, CK => CLK, RN => 
                           n3122, Q => REGISTERS_40_0_port, QN => n_1827);
   REGISTERS_reg_39_31_inst : DFFR_X1 port map( D => n7565, CK => CLK, RN => 
                           n3128, Q => REGISTERS_39_31_port, QN => n_1828);
   REGISTERS_reg_39_30_inst : DFFR_X1 port map( D => n7566, CK => CLK, RN => 
                           n3128, Q => REGISTERS_39_30_port, QN => n_1829);
   REGISTERS_reg_39_29_inst : DFFR_X1 port map( D => n7567, CK => CLK, RN => 
                           n3128, Q => REGISTERS_39_29_port, QN => n_1830);
   REGISTERS_reg_39_28_inst : DFFR_X1 port map( D => n7568, CK => CLK, RN => 
                           n3128, Q => REGISTERS_39_28_port, QN => n_1831);
   REGISTERS_reg_39_27_inst : DFFR_X1 port map( D => n7569, CK => CLK, RN => 
                           n3127, Q => REGISTERS_39_27_port, QN => n_1832);
   REGISTERS_reg_39_26_inst : DFFR_X1 port map( D => n7570, CK => CLK, RN => 
                           n3127, Q => REGISTERS_39_26_port, QN => n_1833);
   REGISTERS_reg_39_25_inst : DFFR_X1 port map( D => n7571, CK => CLK, RN => 
                           n3127, Q => REGISTERS_39_25_port, QN => n_1834);
   REGISTERS_reg_39_24_inst : DFFR_X1 port map( D => n7572, CK => CLK, RN => 
                           n3127, Q => REGISTERS_39_24_port, QN => n_1835);
   REGISTERS_reg_39_23_inst : DFFR_X1 port map( D => n7573, CK => CLK, RN => 
                           n3127, Q => REGISTERS_39_23_port, QN => n_1836);
   REGISTERS_reg_39_22_inst : DFFR_X1 port map( D => n7574, CK => CLK, RN => 
                           n3127, Q => REGISTERS_39_22_port, QN => n_1837);
   REGISTERS_reg_39_21_inst : DFFR_X1 port map( D => n7575, CK => CLK, RN => 
                           n3127, Q => REGISTERS_39_21_port, QN => n_1838);
   REGISTERS_reg_39_20_inst : DFFR_X1 port map( D => n7576, CK => CLK, RN => 
                           n3127, Q => REGISTERS_39_20_port, QN => n_1839);
   REGISTERS_reg_39_19_inst : DFFR_X1 port map( D => n7577, CK => CLK, RN => 
                           n3127, Q => REGISTERS_39_19_port, QN => n_1840);
   REGISTERS_reg_39_18_inst : DFFR_X1 port map( D => n7578, CK => CLK, RN => 
                           n3127, Q => REGISTERS_39_18_port, QN => n_1841);
   REGISTERS_reg_39_17_inst : DFFR_X1 port map( D => n7579, CK => CLK, RN => 
                           n3127, Q => REGISTERS_39_17_port, QN => n_1842);
   REGISTERS_reg_39_16_inst : DFFR_X1 port map( D => n7580, CK => CLK, RN => 
                           n3127, Q => REGISTERS_39_16_port, QN => n_1843);
   REGISTERS_reg_39_15_inst : DFFR_X1 port map( D => n7581, CK => CLK, RN => 
                           n3126, Q => REGISTERS_39_15_port, QN => n_1844);
   REGISTERS_reg_39_14_inst : DFFR_X1 port map( D => n7582, CK => CLK, RN => 
                           n3126, Q => REGISTERS_39_14_port, QN => n_1845);
   REGISTERS_reg_39_13_inst : DFFR_X1 port map( D => n7583, CK => CLK, RN => 
                           n3126, Q => REGISTERS_39_13_port, QN => n_1846);
   REGISTERS_reg_39_12_inst : DFFR_X1 port map( D => n7584, CK => CLK, RN => 
                           n3126, Q => REGISTERS_39_12_port, QN => n_1847);
   REGISTERS_reg_39_11_inst : DFFR_X1 port map( D => n7585, CK => CLK, RN => 
                           n3126, Q => REGISTERS_39_11_port, QN => n_1848);
   REGISTERS_reg_39_10_inst : DFFR_X1 port map( D => n7586, CK => CLK, RN => 
                           n3126, Q => REGISTERS_39_10_port, QN => n_1849);
   REGISTERS_reg_39_9_inst : DFFR_X1 port map( D => n7587, CK => CLK, RN => 
                           n3126, Q => REGISTERS_39_9_port, QN => n_1850);
   REGISTERS_reg_39_8_inst : DFFR_X1 port map( D => n7588, CK => CLK, RN => 
                           n3126, Q => REGISTERS_39_8_port, QN => n_1851);
   REGISTERS_reg_39_7_inst : DFFR_X1 port map( D => n7589, CK => CLK, RN => 
                           n3126, Q => REGISTERS_39_7_port, QN => n_1852);
   REGISTERS_reg_39_6_inst : DFFR_X1 port map( D => n7590, CK => CLK, RN => 
                           n3126, Q => REGISTERS_39_6_port, QN => n_1853);
   REGISTERS_reg_39_5_inst : DFFR_X1 port map( D => n7591, CK => CLK, RN => 
                           n3126, Q => REGISTERS_39_5_port, QN => n_1854);
   REGISTERS_reg_39_4_inst : DFFR_X1 port map( D => n7592, CK => CLK, RN => 
                           n3126, Q => REGISTERS_39_4_port, QN => n_1855);
   REGISTERS_reg_39_3_inst : DFFR_X1 port map( D => n7593, CK => CLK, RN => 
                           n3124, Q => REGISTERS_39_3_port, QN => n_1856);
   REGISTERS_reg_39_2_inst : DFFR_X1 port map( D => n7594, CK => CLK, RN => 
                           n3124, Q => REGISTERS_39_2_port, QN => n_1857);
   REGISTERS_reg_39_1_inst : DFFR_X1 port map( D => n7595, CK => CLK, RN => 
                           n3124, Q => REGISTERS_39_1_port, QN => n_1858);
   REGISTERS_reg_39_0_inst : DFFR_X1 port map( D => n7596, CK => CLK, RN => 
                           n3124, Q => REGISTERS_39_0_port, QN => n_1859);
   REGISTERS_reg_38_31_inst : DFFR_X1 port map( D => n7533, CK => CLK, RN => 
                           n3131, Q => REGISTERS_38_31_port, QN => n_1860);
   REGISTERS_reg_38_30_inst : DFFR_X1 port map( D => n7534, CK => CLK, RN => 
                           n3131, Q => REGISTERS_38_30_port, QN => n_1861);
   REGISTERS_reg_38_29_inst : DFFR_X1 port map( D => n7535, CK => CLK, RN => 
                           n3131, Q => REGISTERS_38_29_port, QN => n_1862);
   REGISTERS_reg_38_28_inst : DFFR_X1 port map( D => n7536, CK => CLK, RN => 
                           n3131, Q => REGISTERS_38_28_port, QN => n_1863);
   REGISTERS_reg_38_27_inst : DFFR_X1 port map( D => n7537, CK => CLK, RN => 
                           n3131, Q => REGISTERS_38_27_port, QN => n_1864);
   REGISTERS_reg_38_26_inst : DFFR_X1 port map( D => n7538, CK => CLK, RN => 
                           n3131, Q => REGISTERS_38_26_port, QN => n_1865);
   REGISTERS_reg_38_25_inst : DFFR_X1 port map( D => n7539, CK => CLK, RN => 
                           n3131, Q => REGISTERS_38_25_port, QN => n_1866);
   REGISTERS_reg_38_24_inst : DFFR_X1 port map( D => n7540, CK => CLK, RN => 
                           n3131, Q => REGISTERS_38_24_port, QN => n_1867);
   REGISTERS_reg_38_23_inst : DFFR_X1 port map( D => n7541, CK => CLK, RN => 
                           n3131, Q => REGISTERS_38_23_port, QN => n_1868);
   REGISTERS_reg_38_22_inst : DFFR_X1 port map( D => n7542, CK => CLK, RN => 
                           n3131, Q => REGISTERS_38_22_port, QN => n_1869);
   REGISTERS_reg_38_21_inst : DFFR_X1 port map( D => n7543, CK => CLK, RN => 
                           n3131, Q => REGISTERS_38_21_port, QN => n_1870);
   REGISTERS_reg_38_20_inst : DFFR_X1 port map( D => n7544, CK => CLK, RN => 
                           n3131, Q => REGISTERS_38_20_port, QN => n_1871);
   REGISTERS_reg_38_19_inst : DFFR_X1 port map( D => n7545, CK => CLK, RN => 
                           n3130, Q => REGISTERS_38_19_port, QN => n_1872);
   REGISTERS_reg_38_18_inst : DFFR_X1 port map( D => n7546, CK => CLK, RN => 
                           n3130, Q => REGISTERS_38_18_port, QN => n_1873);
   REGISTERS_reg_38_17_inst : DFFR_X1 port map( D => n7547, CK => CLK, RN => 
                           n3130, Q => REGISTERS_38_17_port, QN => n_1874);
   REGISTERS_reg_38_16_inst : DFFR_X1 port map( D => n7548, CK => CLK, RN => 
                           n3130, Q => REGISTERS_38_16_port, QN => n_1875);
   REGISTERS_reg_38_15_inst : DFFR_X1 port map( D => n7549, CK => CLK, RN => 
                           n3130, Q => REGISTERS_38_15_port, QN => n_1876);
   REGISTERS_reg_38_14_inst : DFFR_X1 port map( D => n7550, CK => CLK, RN => 
                           n3130, Q => REGISTERS_38_14_port, QN => n_1877);
   REGISTERS_reg_38_13_inst : DFFR_X1 port map( D => n7551, CK => CLK, RN => 
                           n3130, Q => REGISTERS_38_13_port, QN => n_1878);
   REGISTERS_reg_38_12_inst : DFFR_X1 port map( D => n7552, CK => CLK, RN => 
                           n3130, Q => REGISTERS_38_12_port, QN => n_1879);
   REGISTERS_reg_38_11_inst : DFFR_X1 port map( D => n7553, CK => CLK, RN => 
                           n3130, Q => REGISTERS_38_11_port, QN => n_1880);
   REGISTERS_reg_38_10_inst : DFFR_X1 port map( D => n7554, CK => CLK, RN => 
                           n3130, Q => REGISTERS_38_10_port, QN => n_1881);
   REGISTERS_reg_38_9_inst : DFFR_X1 port map( D => n7555, CK => CLK, RN => 
                           n3130, Q => REGISTERS_38_9_port, QN => n_1882);
   REGISTERS_reg_38_8_inst : DFFR_X1 port map( D => n7556, CK => CLK, RN => 
                           n3130, Q => REGISTERS_38_8_port, QN => n_1883);
   REGISTERS_reg_38_7_inst : DFFR_X1 port map( D => n7557, CK => CLK, RN => 
                           n3128, Q => REGISTERS_38_7_port, QN => n_1884);
   REGISTERS_reg_38_6_inst : DFFR_X1 port map( D => n7558, CK => CLK, RN => 
                           n3128, Q => REGISTERS_38_6_port, QN => n_1885);
   REGISTERS_reg_38_5_inst : DFFR_X1 port map( D => n7559, CK => CLK, RN => 
                           n3128, Q => REGISTERS_38_5_port, QN => n_1886);
   REGISTERS_reg_38_4_inst : DFFR_X1 port map( D => n7560, CK => CLK, RN => 
                           n3128, Q => REGISTERS_38_4_port, QN => n_1887);
   REGISTERS_reg_38_3_inst : DFFR_X1 port map( D => n7561, CK => CLK, RN => 
                           n3128, Q => REGISTERS_38_3_port, QN => n_1888);
   REGISTERS_reg_38_2_inst : DFFR_X1 port map( D => n7562, CK => CLK, RN => 
                           n3128, Q => REGISTERS_38_2_port, QN => n_1889);
   REGISTERS_reg_38_1_inst : DFFR_X1 port map( D => n7563, CK => CLK, RN => 
                           n3128, Q => REGISTERS_38_1_port, QN => n_1890);
   REGISTERS_reg_38_0_inst : DFFR_X1 port map( D => n7564, CK => CLK, RN => 
                           n3128, Q => REGISTERS_38_0_port, QN => n_1891);
   REGISTERS_reg_34_31_inst : DFFR_X1 port map( D => n7405, CK => CLK, RN => 
                           n3146, Q => REGISTERS_34_31_port, QN => n_1892);
   REGISTERS_reg_34_30_inst : DFFR_X1 port map( D => n7406, CK => CLK, RN => 
                           n3146, Q => REGISTERS_34_30_port, QN => n_1893);
   REGISTERS_reg_34_29_inst : DFFR_X1 port map( D => n7407, CK => CLK, RN => 
                           n3146, Q => REGISTERS_34_29_port, QN => n_1894);
   REGISTERS_reg_34_28_inst : DFFR_X1 port map( D => n7408, CK => CLK, RN => 
                           n3146, Q => REGISTERS_34_28_port, QN => n_1895);
   REGISTERS_reg_34_27_inst : DFFR_X1 port map( D => n7409, CK => CLK, RN => 
                           n3146, Q => REGISTERS_34_27_port, QN => n_1896);
   REGISTERS_reg_34_26_inst : DFFR_X1 port map( D => n7410, CK => CLK, RN => 
                           n3146, Q => REGISTERS_34_26_port, QN => n_1897);
   REGISTERS_reg_34_25_inst : DFFR_X1 port map( D => n7411, CK => CLK, RN => 
                           n3146, Q => REGISTERS_34_25_port, QN => n_1898);
   REGISTERS_reg_34_24_inst : DFFR_X1 port map( D => n7412, CK => CLK, RN => 
                           n3146, Q => REGISTERS_34_24_port, QN => n_1899);
   REGISTERS_reg_34_23_inst : DFFR_X1 port map( D => n7413, CK => CLK, RN => 
                           n3144, Q => REGISTERS_34_23_port, QN => n_1900);
   REGISTERS_reg_34_22_inst : DFFR_X1 port map( D => n7414, CK => CLK, RN => 
                           n3144, Q => REGISTERS_34_22_port, QN => n_1901);
   REGISTERS_reg_34_21_inst : DFFR_X1 port map( D => n7415, CK => CLK, RN => 
                           n3144, Q => REGISTERS_34_21_port, QN => n_1902);
   REGISTERS_reg_34_20_inst : DFFR_X1 port map( D => n7416, CK => CLK, RN => 
                           n3144, Q => REGISTERS_34_20_port, QN => n_1903);
   REGISTERS_reg_34_19_inst : DFFR_X1 port map( D => n7417, CK => CLK, RN => 
                           n3144, Q => REGISTERS_34_19_port, QN => n_1904);
   REGISTERS_reg_34_18_inst : DFFR_X1 port map( D => n7418, CK => CLK, RN => 
                           n3144, Q => REGISTERS_34_18_port, QN => n_1905);
   REGISTERS_reg_34_17_inst : DFFR_X1 port map( D => n7419, CK => CLK, RN => 
                           n3144, Q => REGISTERS_34_17_port, QN => n_1906);
   REGISTERS_reg_34_16_inst : DFFR_X1 port map( D => n7420, CK => CLK, RN => 
                           n3144, Q => REGISTERS_34_16_port, QN => n_1907);
   REGISTERS_reg_34_15_inst : DFFR_X1 port map( D => n7421, CK => CLK, RN => 
                           n3144, Q => REGISTERS_34_15_port, QN => n_1908);
   REGISTERS_reg_34_14_inst : DFFR_X1 port map( D => n7422, CK => CLK, RN => 
                           n3144, Q => REGISTERS_34_14_port, QN => n_1909);
   REGISTERS_reg_34_13_inst : DFFR_X1 port map( D => n7423, CK => CLK, RN => 
                           n3144, Q => REGISTERS_34_13_port, QN => n_1910);
   REGISTERS_reg_34_12_inst : DFFR_X1 port map( D => n7424, CK => CLK, RN => 
                           n3144, Q => REGISTERS_34_12_port, QN => n_1911);
   REGISTERS_reg_34_11_inst : DFFR_X1 port map( D => n7425, CK => CLK, RN => 
                           n3143, Q => REGISTERS_34_11_port, QN => n_1912);
   REGISTERS_reg_34_10_inst : DFFR_X1 port map( D => n7426, CK => CLK, RN => 
                           n3143, Q => REGISTERS_34_10_port, QN => n_1913);
   REGISTERS_reg_34_9_inst : DFFR_X1 port map( D => n7427, CK => CLK, RN => 
                           n3143, Q => REGISTERS_34_9_port, QN => n_1914);
   REGISTERS_reg_34_8_inst : DFFR_X1 port map( D => n7428, CK => CLK, RN => 
                           n3143, Q => REGISTERS_34_8_port, QN => n_1915);
   REGISTERS_reg_34_7_inst : DFFR_X1 port map( D => n7429, CK => CLK, RN => 
                           n3143, Q => REGISTERS_34_7_port, QN => n_1916);
   REGISTERS_reg_34_6_inst : DFFR_X1 port map( D => n7430, CK => CLK, RN => 
                           n3143, Q => REGISTERS_34_6_port, QN => n_1917);
   REGISTERS_reg_34_5_inst : DFFR_X1 port map( D => n7431, CK => CLK, RN => 
                           n3143, Q => REGISTERS_34_5_port, QN => n_1918);
   REGISTERS_reg_34_4_inst : DFFR_X1 port map( D => n7432, CK => CLK, RN => 
                           n3143, Q => REGISTERS_34_4_port, QN => n_1919);
   REGISTERS_reg_34_3_inst : DFFR_X1 port map( D => n7433, CK => CLK, RN => 
                           n3143, Q => REGISTERS_34_3_port, QN => n_1920);
   REGISTERS_reg_34_2_inst : DFFR_X1 port map( D => n7434, CK => CLK, RN => 
                           n3143, Q => REGISTERS_34_2_port, QN => n_1921);
   REGISTERS_reg_34_1_inst : DFFR_X1 port map( D => n7435, CK => CLK, RN => 
                           n3143, Q => REGISTERS_34_1_port, QN => n_1922);
   REGISTERS_reg_34_0_inst : DFFR_X1 port map( D => n7436, CK => CLK, RN => 
                           n3143, Q => REGISTERS_34_0_port, QN => n_1923);
   REGISTERS_reg_33_31_inst : DFFR_X1 port map( D => n7373, CK => CLK, RN => 
                           n3150, Q => REGISTERS_33_31_port, QN => n_1924);
   REGISTERS_reg_33_30_inst : DFFR_X1 port map( D => n7374, CK => CLK, RN => 
                           n3150, Q => REGISTERS_33_30_port, QN => n_1925);
   REGISTERS_reg_33_29_inst : DFFR_X1 port map( D => n7375, CK => CLK, RN => 
                           n3150, Q => REGISTERS_33_29_port, QN => n_1926);
   REGISTERS_reg_33_28_inst : DFFR_X1 port map( D => n7376, CK => CLK, RN => 
                           n3150, Q => REGISTERS_33_28_port, QN => n_1927);
   REGISTERS_reg_33_27_inst : DFFR_X1 port map( D => n7377, CK => CLK, RN => 
                           n3148, Q => REGISTERS_33_27_port, QN => n_1928);
   REGISTERS_reg_33_26_inst : DFFR_X1 port map( D => n7378, CK => CLK, RN => 
                           n3148, Q => REGISTERS_33_26_port, QN => n_1929);
   REGISTERS_reg_33_25_inst : DFFR_X1 port map( D => n7379, CK => CLK, RN => 
                           n3148, Q => REGISTERS_33_25_port, QN => n_1930);
   REGISTERS_reg_33_24_inst : DFFR_X1 port map( D => n7380, CK => CLK, RN => 
                           n3148, Q => REGISTERS_33_24_port, QN => n_1931);
   REGISTERS_reg_33_23_inst : DFFR_X1 port map( D => n7381, CK => CLK, RN => 
                           n3148, Q => REGISTERS_33_23_port, QN => n_1932);
   REGISTERS_reg_33_22_inst : DFFR_X1 port map( D => n7382, CK => CLK, RN => 
                           n3148, Q => REGISTERS_33_22_port, QN => n_1933);
   REGISTERS_reg_33_21_inst : DFFR_X1 port map( D => n7383, CK => CLK, RN => 
                           n3148, Q => REGISTERS_33_21_port, QN => n_1934);
   REGISTERS_reg_33_20_inst : DFFR_X1 port map( D => n7384, CK => CLK, RN => 
                           n3148, Q => REGISTERS_33_20_port, QN => n_1935);
   REGISTERS_reg_33_19_inst : DFFR_X1 port map( D => n7385, CK => CLK, RN => 
                           n3148, Q => REGISTERS_33_19_port, QN => n_1936);
   REGISTERS_reg_33_18_inst : DFFR_X1 port map( D => n7386, CK => CLK, RN => 
                           n3148, Q => REGISTERS_33_18_port, QN => n_1937);
   REGISTERS_reg_33_17_inst : DFFR_X1 port map( D => n7387, CK => CLK, RN => 
                           n3148, Q => REGISTERS_33_17_port, QN => n_1938);
   REGISTERS_reg_33_16_inst : DFFR_X1 port map( D => n7388, CK => CLK, RN => 
                           n3148, Q => REGISTERS_33_16_port, QN => n_1939);
   REGISTERS_reg_33_15_inst : DFFR_X1 port map( D => n7389, CK => CLK, RN => 
                           n3147, Q => REGISTERS_33_15_port, QN => n_1940);
   REGISTERS_reg_33_14_inst : DFFR_X1 port map( D => n7390, CK => CLK, RN => 
                           n3147, Q => REGISTERS_33_14_port, QN => n_1941);
   REGISTERS_reg_33_13_inst : DFFR_X1 port map( D => n7391, CK => CLK, RN => 
                           n3147, Q => REGISTERS_33_13_port, QN => n_1942);
   REGISTERS_reg_33_12_inst : DFFR_X1 port map( D => n7392, CK => CLK, RN => 
                           n3147, Q => REGISTERS_33_12_port, QN => n_1943);
   REGISTERS_reg_33_11_inst : DFFR_X1 port map( D => n7393, CK => CLK, RN => 
                           n3147, Q => REGISTERS_33_11_port, QN => n_1944);
   REGISTERS_reg_33_10_inst : DFFR_X1 port map( D => n7394, CK => CLK, RN => 
                           n3147, Q => REGISTERS_33_10_port, QN => n_1945);
   REGISTERS_reg_33_9_inst : DFFR_X1 port map( D => n7395, CK => CLK, RN => 
                           n3147, Q => REGISTERS_33_9_port, QN => n_1946);
   REGISTERS_reg_33_8_inst : DFFR_X1 port map( D => n7396, CK => CLK, RN => 
                           n3147, Q => REGISTERS_33_8_port, QN => n_1947);
   REGISTERS_reg_33_7_inst : DFFR_X1 port map( D => n7397, CK => CLK, RN => 
                           n3147, Q => REGISTERS_33_7_port, QN => n_1948);
   REGISTERS_reg_33_6_inst : DFFR_X1 port map( D => n7398, CK => CLK, RN => 
                           n3147, Q => REGISTERS_33_6_port, QN => n_1949);
   REGISTERS_reg_33_5_inst : DFFR_X1 port map( D => n7399, CK => CLK, RN => 
                           n3147, Q => REGISTERS_33_5_port, QN => n_1950);
   REGISTERS_reg_33_4_inst : DFFR_X1 port map( D => n7400, CK => CLK, RN => 
                           n3147, Q => REGISTERS_33_4_port, QN => n_1951);
   REGISTERS_reg_33_3_inst : DFFR_X1 port map( D => n7401, CK => CLK, RN => 
                           n3146, Q => REGISTERS_33_3_port, QN => n_1952);
   REGISTERS_reg_33_2_inst : DFFR_X1 port map( D => n7402, CK => CLK, RN => 
                           n3146, Q => REGISTERS_33_2_port, QN => n_1953);
   REGISTERS_reg_33_1_inst : DFFR_X1 port map( D => n7403, CK => CLK, RN => 
                           n3146, Q => REGISTERS_33_1_port, QN => n_1954);
   REGISTERS_reg_33_0_inst : DFFR_X1 port map( D => n7404, CK => CLK, RN => 
                           n3146, Q => REGISTERS_33_0_port, QN => n_1955);
   REGISTERS_reg_21_31_inst : DFFR_X1 port map( D => n6989, CK => CLK, RN => 
                           n3193, Q => REGISTERS_21_31_port, QN => n_1956);
   REGISTERS_reg_21_30_inst : DFFR_X1 port map( D => n6990, CK => CLK, RN => 
                           n3193, Q => REGISTERS_21_30_port, QN => n_1957);
   REGISTERS_reg_21_29_inst : DFFR_X1 port map( D => n6991, CK => CLK, RN => 
                           n3193, Q => REGISTERS_21_29_port, QN => n_1958);
   REGISTERS_reg_21_28_inst : DFFR_X1 port map( D => n6992, CK => CLK, RN => 
                           n3193, Q => REGISTERS_21_28_port, QN => n_1959);
   REGISTERS_reg_21_27_inst : DFFR_X1 port map( D => n6993, CK => CLK, RN => 
                           n3192, Q => REGISTERS_21_27_port, QN => n_1960);
   REGISTERS_reg_21_26_inst : DFFR_X1 port map( D => n6994, CK => CLK, RN => 
                           n3192, Q => REGISTERS_21_26_port, QN => n_1961);
   REGISTERS_reg_21_25_inst : DFFR_X1 port map( D => n6995, CK => CLK, RN => 
                           n3192, Q => REGISTERS_21_25_port, QN => n_1962);
   REGISTERS_reg_21_24_inst : DFFR_X1 port map( D => n6996, CK => CLK, RN => 
                           n3192, Q => REGISTERS_21_24_port, QN => n_1963);
   REGISTERS_reg_21_23_inst : DFFR_X1 port map( D => n6997, CK => CLK, RN => 
                           n3192, Q => REGISTERS_21_23_port, QN => n_1964);
   REGISTERS_reg_21_22_inst : DFFR_X1 port map( D => n6998, CK => CLK, RN => 
                           n3192, Q => REGISTERS_21_22_port, QN => n_1965);
   REGISTERS_reg_21_21_inst : DFFR_X1 port map( D => n6999, CK => CLK, RN => 
                           n3192, Q => REGISTERS_21_21_port, QN => n_1966);
   REGISTERS_reg_21_20_inst : DFFR_X1 port map( D => n7000, CK => CLK, RN => 
                           n3192, Q => REGISTERS_21_20_port, QN => n_1967);
   REGISTERS_reg_21_19_inst : DFFR_X1 port map( D => n7001, CK => CLK, RN => 
                           n3192, Q => REGISTERS_21_19_port, QN => n_1968);
   REGISTERS_reg_21_18_inst : DFFR_X1 port map( D => n7002, CK => CLK, RN => 
                           n3192, Q => REGISTERS_21_18_port, QN => n_1969);
   REGISTERS_reg_21_17_inst : DFFR_X1 port map( D => n7003, CK => CLK, RN => 
                           n3192, Q => REGISTERS_21_17_port, QN => n_1970);
   REGISTERS_reg_21_16_inst : DFFR_X1 port map( D => n7004, CK => CLK, RN => 
                           n3192, Q => REGISTERS_21_16_port, QN => n_1971);
   REGISTERS_reg_21_15_inst : DFFR_X1 port map( D => n7005, CK => CLK, RN => 
                           n3191, Q => REGISTERS_21_15_port, QN => n_1972);
   REGISTERS_reg_21_14_inst : DFFR_X1 port map( D => n7006, CK => CLK, RN => 
                           n3191, Q => REGISTERS_21_14_port, QN => n_1973);
   REGISTERS_reg_21_13_inst : DFFR_X1 port map( D => n7007, CK => CLK, RN => 
                           n3191, Q => REGISTERS_21_13_port, QN => n_1974);
   REGISTERS_reg_21_12_inst : DFFR_X1 port map( D => n7008, CK => CLK, RN => 
                           n3191, Q => REGISTERS_21_12_port, QN => n_1975);
   REGISTERS_reg_21_11_inst : DFFR_X1 port map( D => n7009, CK => CLK, RN => 
                           n3191, Q => REGISTERS_21_11_port, QN => n_1976);
   REGISTERS_reg_21_10_inst : DFFR_X1 port map( D => n7010, CK => CLK, RN => 
                           n3191, Q => REGISTERS_21_10_port, QN => n_1977);
   REGISTERS_reg_21_9_inst : DFFR_X1 port map( D => n7011, CK => CLK, RN => 
                           n3191, Q => REGISTERS_21_9_port, QN => n_1978);
   REGISTERS_reg_21_8_inst : DFFR_X1 port map( D => n7012, CK => CLK, RN => 
                           n3191, Q => REGISTERS_21_8_port, QN => n_1979);
   REGISTERS_reg_21_7_inst : DFFR_X1 port map( D => n7013, CK => CLK, RN => 
                           n3191, Q => REGISTERS_21_7_port, QN => n_1980);
   REGISTERS_reg_21_6_inst : DFFR_X1 port map( D => n7014, CK => CLK, RN => 
                           n3191, Q => REGISTERS_21_6_port, QN => n_1981);
   REGISTERS_reg_21_5_inst : DFFR_X1 port map( D => n7015, CK => CLK, RN => 
                           n3191, Q => REGISTERS_21_5_port, QN => n_1982);
   REGISTERS_reg_21_4_inst : DFFR_X1 port map( D => n7016, CK => CLK, RN => 
                           n3191, Q => REGISTERS_21_4_port, QN => n_1983);
   REGISTERS_reg_21_3_inst : DFFR_X1 port map( D => n7017, CK => CLK, RN => 
                           n3189, Q => REGISTERS_21_3_port, QN => n_1984);
   REGISTERS_reg_21_2_inst : DFFR_X1 port map( D => n7018, CK => CLK, RN => 
                           n3189, Q => REGISTERS_21_2_port, QN => n_1985);
   REGISTERS_reg_21_1_inst : DFFR_X1 port map( D => n7019, CK => CLK, RN => 
                           n3189, Q => REGISTERS_21_1_port, QN => n_1986);
   REGISTERS_reg_21_0_inst : DFFR_X1 port map( D => n7020, CK => CLK, RN => 
                           n3189, Q => REGISTERS_21_0_port, QN => n_1987);
   REGISTERS_reg_20_31_inst : DFFR_X1 port map( D => n6957, CK => CLK, RN => 
                           n3196, Q => REGISTERS_20_31_port, QN => n_1988);
   REGISTERS_reg_20_30_inst : DFFR_X1 port map( D => n6958, CK => CLK, RN => 
                           n3196, Q => REGISTERS_20_30_port, QN => n_1989);
   REGISTERS_reg_20_29_inst : DFFR_X1 port map( D => n6959, CK => CLK, RN => 
                           n3196, Q => REGISTERS_20_29_port, QN => n_1990);
   REGISTERS_reg_20_28_inst : DFFR_X1 port map( D => n6960, CK => CLK, RN => 
                           n3196, Q => REGISTERS_20_28_port, QN => n_1991);
   REGISTERS_reg_20_27_inst : DFFR_X1 port map( D => n6961, CK => CLK, RN => 
                           n3196, Q => REGISTERS_20_27_port, QN => n_1992);
   REGISTERS_reg_20_26_inst : DFFR_X1 port map( D => n6962, CK => CLK, RN => 
                           n3196, Q => REGISTERS_20_26_port, QN => n_1993);
   REGISTERS_reg_20_25_inst : DFFR_X1 port map( D => n6963, CK => CLK, RN => 
                           n3196, Q => REGISTERS_20_25_port, QN => n_1994);
   REGISTERS_reg_20_24_inst : DFFR_X1 port map( D => n6964, CK => CLK, RN => 
                           n3196, Q => REGISTERS_20_24_port, QN => n_1995);
   REGISTERS_reg_20_23_inst : DFFR_X1 port map( D => n6965, CK => CLK, RN => 
                           n3196, Q => REGISTERS_20_23_port, QN => n_1996);
   REGISTERS_reg_20_22_inst : DFFR_X1 port map( D => n6966, CK => CLK, RN => 
                           n3196, Q => REGISTERS_20_22_port, QN => n_1997);
   REGISTERS_reg_20_21_inst : DFFR_X1 port map( D => n6967, CK => CLK, RN => 
                           n3196, Q => REGISTERS_20_21_port, QN => n_1998);
   REGISTERS_reg_20_20_inst : DFFR_X1 port map( D => n6968, CK => CLK, RN => 
                           n3196, Q => REGISTERS_20_20_port, QN => n_1999);
   REGISTERS_reg_20_19_inst : DFFR_X1 port map( D => n6969, CK => CLK, RN => 
                           n3195, Q => REGISTERS_20_19_port, QN => n_2000);
   REGISTERS_reg_20_18_inst : DFFR_X1 port map( D => n6970, CK => CLK, RN => 
                           n3195, Q => REGISTERS_20_18_port, QN => n_2001);
   REGISTERS_reg_20_17_inst : DFFR_X1 port map( D => n6971, CK => CLK, RN => 
                           n3195, Q => REGISTERS_20_17_port, QN => n_2002);
   REGISTERS_reg_20_16_inst : DFFR_X1 port map( D => n6972, CK => CLK, RN => 
                           n3195, Q => REGISTERS_20_16_port, QN => n_2003);
   REGISTERS_reg_20_15_inst : DFFR_X1 port map( D => n6973, CK => CLK, RN => 
                           n3195, Q => REGISTERS_20_15_port, QN => n_2004);
   REGISTERS_reg_20_14_inst : DFFR_X1 port map( D => n6974, CK => CLK, RN => 
                           n3195, Q => REGISTERS_20_14_port, QN => n_2005);
   REGISTERS_reg_20_13_inst : DFFR_X1 port map( D => n6975, CK => CLK, RN => 
                           n3195, Q => REGISTERS_20_13_port, QN => n_2006);
   REGISTERS_reg_20_12_inst : DFFR_X1 port map( D => n6976, CK => CLK, RN => 
                           n3195, Q => REGISTERS_20_12_port, QN => n_2007);
   REGISTERS_reg_20_11_inst : DFFR_X1 port map( D => n6977, CK => CLK, RN => 
                           n3195, Q => REGISTERS_20_11_port, QN => n_2008);
   REGISTERS_reg_20_10_inst : DFFR_X1 port map( D => n6978, CK => CLK, RN => 
                           n3195, Q => REGISTERS_20_10_port, QN => n_2009);
   REGISTERS_reg_20_9_inst : DFFR_X1 port map( D => n6979, CK => CLK, RN => 
                           n3195, Q => REGISTERS_20_9_port, QN => n_2010);
   REGISTERS_reg_20_8_inst : DFFR_X1 port map( D => n6980, CK => CLK, RN => 
                           n3195, Q => REGISTERS_20_8_port, QN => n_2011);
   REGISTERS_reg_20_7_inst : DFFR_X1 port map( D => n6981, CK => CLK, RN => 
                           n3193, Q => REGISTERS_20_7_port, QN => n_2012);
   REGISTERS_reg_20_6_inst : DFFR_X1 port map( D => n6982, CK => CLK, RN => 
                           n3193, Q => REGISTERS_20_6_port, QN => n_2013);
   REGISTERS_reg_20_5_inst : DFFR_X1 port map( D => n6983, CK => CLK, RN => 
                           n3193, Q => REGISTERS_20_5_port, QN => n_2014);
   REGISTERS_reg_20_4_inst : DFFR_X1 port map( D => n6984, CK => CLK, RN => 
                           n3193, Q => REGISTERS_20_4_port, QN => n_2015);
   REGISTERS_reg_20_3_inst : DFFR_X1 port map( D => n6985, CK => CLK, RN => 
                           n3193, Q => REGISTERS_20_3_port, QN => n_2016);
   REGISTERS_reg_20_2_inst : DFFR_X1 port map( D => n6986, CK => CLK, RN => 
                           n3193, Q => REGISTERS_20_2_port, QN => n_2017);
   REGISTERS_reg_20_1_inst : DFFR_X1 port map( D => n6987, CK => CLK, RN => 
                           n3193, Q => REGISTERS_20_1_port, QN => n_2018);
   REGISTERS_reg_20_0_inst : DFFR_X1 port map( D => n6988, CK => CLK, RN => 
                           n3193, Q => REGISTERS_20_0_port, QN => n_2019);
   REGISTERS_reg_19_31_inst : DFFR_X1 port map( D => n6925, CK => CLK, RN => 
                           n3200, Q => REGISTERS_19_31_port, QN => n_2020);
   REGISTERS_reg_19_30_inst : DFFR_X1 port map( D => n6926, CK => CLK, RN => 
                           n3200, Q => REGISTERS_19_30_port, QN => n_2021);
   REGISTERS_reg_19_29_inst : DFFR_X1 port map( D => n6927, CK => CLK, RN => 
                           n3200, Q => REGISTERS_19_29_port, QN => n_2022);
   REGISTERS_reg_19_28_inst : DFFR_X1 port map( D => n6928, CK => CLK, RN => 
                           n3200, Q => REGISTERS_19_28_port, QN => n_2023);
   REGISTERS_reg_19_27_inst : DFFR_X1 port map( D => n6929, CK => CLK, RN => 
                           n3200, Q => REGISTERS_19_27_port, QN => n_2024);
   REGISTERS_reg_19_26_inst : DFFR_X1 port map( D => n6930, CK => CLK, RN => 
                           n3200, Q => REGISTERS_19_26_port, QN => n_2025);
   REGISTERS_reg_19_25_inst : DFFR_X1 port map( D => n6931, CK => CLK, RN => 
                           n3200, Q => REGISTERS_19_25_port, QN => n_2026);
   REGISTERS_reg_19_24_inst : DFFR_X1 port map( D => n6932, CK => CLK, RN => 
                           n3200, Q => REGISTERS_19_24_port, QN => n_2027);
   REGISTERS_reg_19_23_inst : DFFR_X1 port map( D => n6933, CK => CLK, RN => 
                           n3199, Q => REGISTERS_19_23_port, QN => n_2028);
   REGISTERS_reg_19_22_inst : DFFR_X1 port map( D => n6934, CK => CLK, RN => 
                           n3199, Q => REGISTERS_19_22_port, QN => n_2029);
   REGISTERS_reg_19_21_inst : DFFR_X1 port map( D => n6935, CK => CLK, RN => 
                           n3199, Q => REGISTERS_19_21_port, QN => n_2030);
   REGISTERS_reg_19_20_inst : DFFR_X1 port map( D => n6936, CK => CLK, RN => 
                           n3199, Q => REGISTERS_19_20_port, QN => n_2031);
   REGISTERS_reg_19_19_inst : DFFR_X1 port map( D => n6937, CK => CLK, RN => 
                           n3199, Q => REGISTERS_19_19_port, QN => n_2032);
   REGISTERS_reg_19_18_inst : DFFR_X1 port map( D => n6938, CK => CLK, RN => 
                           n3199, Q => REGISTERS_19_18_port, QN => n_2033);
   REGISTERS_reg_19_17_inst : DFFR_X1 port map( D => n6939, CK => CLK, RN => 
                           n3199, Q => REGISTERS_19_17_port, QN => n_2034);
   REGISTERS_reg_19_16_inst : DFFR_X1 port map( D => n6940, CK => CLK, RN => 
                           n3199, Q => REGISTERS_19_16_port, QN => n_2035);
   REGISTERS_reg_19_15_inst : DFFR_X1 port map( D => n6941, CK => CLK, RN => 
                           n3199, Q => REGISTERS_19_15_port, QN => n_2036);
   REGISTERS_reg_19_14_inst : DFFR_X1 port map( D => n6942, CK => CLK, RN => 
                           n3199, Q => REGISTERS_19_14_port, QN => n_2037);
   REGISTERS_reg_19_13_inst : DFFR_X1 port map( D => n6943, CK => CLK, RN => 
                           n3199, Q => REGISTERS_19_13_port, QN => n_2038);
   REGISTERS_reg_19_12_inst : DFFR_X1 port map( D => n6944, CK => CLK, RN => 
                           n3199, Q => REGISTERS_19_12_port, QN => n_2039);
   REGISTERS_reg_19_11_inst : DFFR_X1 port map( D => n6945, CK => CLK, RN => 
                           n3197, Q => REGISTERS_19_11_port, QN => n_2040);
   REGISTERS_reg_19_10_inst : DFFR_X1 port map( D => n6946, CK => CLK, RN => 
                           n3197, Q => REGISTERS_19_10_port, QN => n_2041);
   REGISTERS_reg_19_9_inst : DFFR_X1 port map( D => n6947, CK => CLK, RN => 
                           n3197, Q => REGISTERS_19_9_port, QN => n_2042);
   REGISTERS_reg_19_8_inst : DFFR_X1 port map( D => n6948, CK => CLK, RN => 
                           n3197, Q => REGISTERS_19_8_port, QN => n_2043);
   REGISTERS_reg_19_7_inst : DFFR_X1 port map( D => n6949, CK => CLK, RN => 
                           n3197, Q => REGISTERS_19_7_port, QN => n_2044);
   REGISTERS_reg_19_6_inst : DFFR_X1 port map( D => n6950, CK => CLK, RN => 
                           n3197, Q => REGISTERS_19_6_port, QN => n_2045);
   REGISTERS_reg_19_5_inst : DFFR_X1 port map( D => n6951, CK => CLK, RN => 
                           n3197, Q => REGISTERS_19_5_port, QN => n_2046);
   REGISTERS_reg_19_4_inst : DFFR_X1 port map( D => n6952, CK => CLK, RN => 
                           n3197, Q => REGISTERS_19_4_port, QN => n_2047);
   REGISTERS_reg_19_3_inst : DFFR_X1 port map( D => n6953, CK => CLK, RN => 
                           n3197, Q => REGISTERS_19_3_port, QN => n_2048);
   REGISTERS_reg_19_2_inst : DFFR_X1 port map( D => n6954, CK => CLK, RN => 
                           n3197, Q => REGISTERS_19_2_port, QN => n_2049);
   REGISTERS_reg_19_1_inst : DFFR_X1 port map( D => n6955, CK => CLK, RN => 
                           n3197, Q => REGISTERS_19_1_port, QN => n_2050);
   REGISTERS_reg_19_0_inst : DFFR_X1 port map( D => n6956, CK => CLK, RN => 
                           n3197, Q => REGISTERS_19_0_port, QN => n_2051);
   REGISTERS_reg_18_31_inst : DFFR_X1 port map( D => n6893, CK => CLK, RN => 
                           n3204, Q => REGISTERS_18_31_port, QN => n_2052);
   REGISTERS_reg_18_30_inst : DFFR_X1 port map( D => n6894, CK => CLK, RN => 
                           n3204, Q => REGISTERS_18_30_port, QN => n_2053);
   REGISTERS_reg_18_29_inst : DFFR_X1 port map( D => n6895, CK => CLK, RN => 
                           n3204, Q => REGISTERS_18_29_port, QN => n_2054);
   REGISTERS_reg_18_28_inst : DFFR_X1 port map( D => n6896, CK => CLK, RN => 
                           n3204, Q => REGISTERS_18_28_port, QN => n_2055);
   REGISTERS_reg_18_27_inst : DFFR_X1 port map( D => n6897, CK => CLK, RN => 
                           n3203, Q => REGISTERS_18_27_port, QN => n_2056);
   REGISTERS_reg_18_26_inst : DFFR_X1 port map( D => n6898, CK => CLK, RN => 
                           n3203, Q => REGISTERS_18_26_port, QN => n_2057);
   REGISTERS_reg_18_25_inst : DFFR_X1 port map( D => n6899, CK => CLK, RN => 
                           n3203, Q => REGISTERS_18_25_port, QN => n_2058);
   REGISTERS_reg_18_24_inst : DFFR_X1 port map( D => n6900, CK => CLK, RN => 
                           n3203, Q => REGISTERS_18_24_port, QN => n_2059);
   REGISTERS_reg_18_23_inst : DFFR_X1 port map( D => n6901, CK => CLK, RN => 
                           n3203, Q => REGISTERS_18_23_port, QN => n_2060);
   REGISTERS_reg_18_22_inst : DFFR_X1 port map( D => n6902, CK => CLK, RN => 
                           n3203, Q => REGISTERS_18_22_port, QN => n_2061);
   REGISTERS_reg_18_21_inst : DFFR_X1 port map( D => n6903, CK => CLK, RN => 
                           n3203, Q => REGISTERS_18_21_port, QN => n_2062);
   REGISTERS_reg_18_20_inst : DFFR_X1 port map( D => n6904, CK => CLK, RN => 
                           n3203, Q => REGISTERS_18_20_port, QN => n_2063);
   REGISTERS_reg_18_19_inst : DFFR_X1 port map( D => n6905, CK => CLK, RN => 
                           n3203, Q => REGISTERS_18_19_port, QN => n_2064);
   REGISTERS_reg_18_18_inst : DFFR_X1 port map( D => n6906, CK => CLK, RN => 
                           n3203, Q => REGISTERS_18_18_port, QN => n_2065);
   REGISTERS_reg_18_17_inst : DFFR_X1 port map( D => n6907, CK => CLK, RN => 
                           n3203, Q => REGISTERS_18_17_port, QN => n_2066);
   REGISTERS_reg_18_16_inst : DFFR_X1 port map( D => n6908, CK => CLK, RN => 
                           n3203, Q => REGISTERS_18_16_port, QN => n_2067);
   REGISTERS_reg_18_15_inst : DFFR_X1 port map( D => n6909, CK => CLK, RN => 
                           n3201, Q => REGISTERS_18_15_port, QN => n_2068);
   REGISTERS_reg_18_14_inst : DFFR_X1 port map( D => n6910, CK => CLK, RN => 
                           n3201, Q => REGISTERS_18_14_port, QN => n_2069);
   REGISTERS_reg_18_13_inst : DFFR_X1 port map( D => n6911, CK => CLK, RN => 
                           n3201, Q => REGISTERS_18_13_port, QN => n_2070);
   REGISTERS_reg_18_12_inst : DFFR_X1 port map( D => n6912, CK => CLK, RN => 
                           n3201, Q => REGISTERS_18_12_port, QN => n_2071);
   REGISTERS_reg_18_11_inst : DFFR_X1 port map( D => n6913, CK => CLK, RN => 
                           n3201, Q => REGISTERS_18_11_port, QN => n_2072);
   REGISTERS_reg_18_10_inst : DFFR_X1 port map( D => n6914, CK => CLK, RN => 
                           n3201, Q => REGISTERS_18_10_port, QN => n_2073);
   REGISTERS_reg_18_9_inst : DFFR_X1 port map( D => n6915, CK => CLK, RN => 
                           n3201, Q => REGISTERS_18_9_port, QN => n_2074);
   REGISTERS_reg_18_8_inst : DFFR_X1 port map( D => n6916, CK => CLK, RN => 
                           n3201, Q => REGISTERS_18_8_port, QN => n_2075);
   REGISTERS_reg_18_7_inst : DFFR_X1 port map( D => n6917, CK => CLK, RN => 
                           n3201, Q => REGISTERS_18_7_port, QN => n_2076);
   REGISTERS_reg_18_6_inst : DFFR_X1 port map( D => n6918, CK => CLK, RN => 
                           n3201, Q => REGISTERS_18_6_port, QN => n_2077);
   REGISTERS_reg_18_5_inst : DFFR_X1 port map( D => n6919, CK => CLK, RN => 
                           n3201, Q => REGISTERS_18_5_port, QN => n_2078);
   REGISTERS_reg_18_4_inst : DFFR_X1 port map( D => n6920, CK => CLK, RN => 
                           n3201, Q => REGISTERS_18_4_port, QN => n_2079);
   REGISTERS_reg_18_3_inst : DFFR_X1 port map( D => n6921, CK => CLK, RN => 
                           n3200, Q => REGISTERS_18_3_port, QN => n_2080);
   REGISTERS_reg_18_2_inst : DFFR_X1 port map( D => n6922, CK => CLK, RN => 
                           n3200, Q => REGISTERS_18_2_port, QN => n_2081);
   REGISTERS_reg_18_1_inst : DFFR_X1 port map( D => n6923, CK => CLK, RN => 
                           n3200, Q => REGISTERS_18_1_port, QN => n_2082);
   REGISTERS_reg_18_0_inst : DFFR_X1 port map( D => n6924, CK => CLK, RN => 
                           n3200, Q => REGISTERS_18_0_port, QN => n_2083);
   REGISTERS_reg_17_31_inst : DFFR_X1 port map( D => n6861, CK => CLK, RN => 
                           n3207, Q => REGISTERS_17_31_port, QN => n_2084);
   REGISTERS_reg_17_30_inst : DFFR_X1 port map( D => n6862, CK => CLK, RN => 
                           n3207, Q => REGISTERS_17_30_port, QN => n_2085);
   REGISTERS_reg_17_29_inst : DFFR_X1 port map( D => n6863, CK => CLK, RN => 
                           n3207, Q => REGISTERS_17_29_port, QN => n_2086);
   REGISTERS_reg_17_28_inst : DFFR_X1 port map( D => n6864, CK => CLK, RN => 
                           n3207, Q => REGISTERS_17_28_port, QN => n_2087);
   REGISTERS_reg_17_27_inst : DFFR_X1 port map( D => n6865, CK => CLK, RN => 
                           n3207, Q => REGISTERS_17_27_port, QN => n_2088);
   REGISTERS_reg_17_26_inst : DFFR_X1 port map( D => n6866, CK => CLK, RN => 
                           n3207, Q => REGISTERS_17_26_port, QN => n_2089);
   REGISTERS_reg_17_25_inst : DFFR_X1 port map( D => n6867, CK => CLK, RN => 
                           n3207, Q => REGISTERS_17_25_port, QN => n_2090);
   REGISTERS_reg_17_24_inst : DFFR_X1 port map( D => n6868, CK => CLK, RN => 
                           n3207, Q => REGISTERS_17_24_port, QN => n_2091);
   REGISTERS_reg_17_23_inst : DFFR_X1 port map( D => n6869, CK => CLK, RN => 
                           n3207, Q => REGISTERS_17_23_port, QN => n_2092);
   REGISTERS_reg_17_22_inst : DFFR_X1 port map( D => n6870, CK => CLK, RN => 
                           n3207, Q => REGISTERS_17_22_port, QN => n_2093);
   REGISTERS_reg_17_21_inst : DFFR_X1 port map( D => n6871, CK => CLK, RN => 
                           n3207, Q => REGISTERS_17_21_port, QN => n_2094);
   REGISTERS_reg_17_20_inst : DFFR_X1 port map( D => n6872, CK => CLK, RN => 
                           n3207, Q => REGISTERS_17_20_port, QN => n_2095);
   REGISTERS_reg_17_19_inst : DFFR_X1 port map( D => n6873, CK => CLK, RN => 
                           n3205, Q => REGISTERS_17_19_port, QN => n_2096);
   REGISTERS_reg_17_18_inst : DFFR_X1 port map( D => n6874, CK => CLK, RN => 
                           n3205, Q => REGISTERS_17_18_port, QN => n_2097);
   REGISTERS_reg_17_17_inst : DFFR_X1 port map( D => n6875, CK => CLK, RN => 
                           n3205, Q => REGISTERS_17_17_port, QN => n_2098);
   REGISTERS_reg_17_16_inst : DFFR_X1 port map( D => n6876, CK => CLK, RN => 
                           n3205, Q => REGISTERS_17_16_port, QN => n_2099);
   REGISTERS_reg_17_15_inst : DFFR_X1 port map( D => n6877, CK => CLK, RN => 
                           n3205, Q => REGISTERS_17_15_port, QN => n_2100);
   REGISTERS_reg_17_14_inst : DFFR_X1 port map( D => n6878, CK => CLK, RN => 
                           n3205, Q => REGISTERS_17_14_port, QN => n_2101);
   REGISTERS_reg_17_13_inst : DFFR_X1 port map( D => n6879, CK => CLK, RN => 
                           n3205, Q => REGISTERS_17_13_port, QN => n_2102);
   REGISTERS_reg_17_12_inst : DFFR_X1 port map( D => n6880, CK => CLK, RN => 
                           n3205, Q => REGISTERS_17_12_port, QN => n_2103);
   REGISTERS_reg_17_11_inst : DFFR_X1 port map( D => n6881, CK => CLK, RN => 
                           n3205, Q => REGISTERS_17_11_port, QN => n_2104);
   REGISTERS_reg_17_10_inst : DFFR_X1 port map( D => n6882, CK => CLK, RN => 
                           n3205, Q => REGISTERS_17_10_port, QN => n_2105);
   REGISTERS_reg_17_9_inst : DFFR_X1 port map( D => n6883, CK => CLK, RN => 
                           n3205, Q => REGISTERS_17_9_port, QN => n_2106);
   REGISTERS_reg_17_8_inst : DFFR_X1 port map( D => n6884, CK => CLK, RN => 
                           n3205, Q => REGISTERS_17_8_port, QN => n_2107);
   REGISTERS_reg_17_7_inst : DFFR_X1 port map( D => n6885, CK => CLK, RN => 
                           n3204, Q => REGISTERS_17_7_port, QN => n_2108);
   REGISTERS_reg_17_6_inst : DFFR_X1 port map( D => n6886, CK => CLK, RN => 
                           n3204, Q => REGISTERS_17_6_port, QN => n_2109);
   REGISTERS_reg_17_5_inst : DFFR_X1 port map( D => n6887, CK => CLK, RN => 
                           n3204, Q => REGISTERS_17_5_port, QN => n_2110);
   REGISTERS_reg_17_4_inst : DFFR_X1 port map( D => n6888, CK => CLK, RN => 
                           n3204, Q => REGISTERS_17_4_port, QN => n_2111);
   REGISTERS_reg_17_3_inst : DFFR_X1 port map( D => n6889, CK => CLK, RN => 
                           n3204, Q => REGISTERS_17_3_port, QN => n_2112);
   REGISTERS_reg_17_2_inst : DFFR_X1 port map( D => n6890, CK => CLK, RN => 
                           n3204, Q => REGISTERS_17_2_port, QN => n_2113);
   REGISTERS_reg_17_1_inst : DFFR_X1 port map( D => n6891, CK => CLK, RN => 
                           n3204, Q => REGISTERS_17_1_port, QN => n_2114);
   REGISTERS_reg_17_0_inst : DFFR_X1 port map( D => n6892, CK => CLK, RN => 
                           n3204, Q => REGISTERS_17_0_port, QN => n_2115);
   REGISTERS_reg_16_31_inst : DFFR_X1 port map( D => n6829, CK => CLK, RN => 
                           n3211, Q => REGISTERS_16_31_port, QN => n_2116);
   REGISTERS_reg_16_30_inst : DFFR_X1 port map( D => n6830, CK => CLK, RN => 
                           n3211, Q => REGISTERS_16_30_port, QN => n_2117);
   REGISTERS_reg_16_29_inst : DFFR_X1 port map( D => n6831, CK => CLK, RN => 
                           n3211, Q => REGISTERS_16_29_port, QN => n_2118);
   REGISTERS_reg_16_28_inst : DFFR_X1 port map( D => n6832, CK => CLK, RN => 
                           n3211, Q => REGISTERS_16_28_port, QN => n_2119);
   REGISTERS_reg_16_27_inst : DFFR_X1 port map( D => n6833, CK => CLK, RN => 
                           n3211, Q => REGISTERS_16_27_port, QN => n_2120);
   REGISTERS_reg_16_26_inst : DFFR_X1 port map( D => n6834, CK => CLK, RN => 
                           n3211, Q => REGISTERS_16_26_port, QN => n_2121);
   REGISTERS_reg_16_25_inst : DFFR_X1 port map( D => n6835, CK => CLK, RN => 
                           n3211, Q => REGISTERS_16_25_port, QN => n_2122);
   REGISTERS_reg_16_24_inst : DFFR_X1 port map( D => n6836, CK => CLK, RN => 
                           n3211, Q => REGISTERS_16_24_port, QN => n_2123);
   REGISTERS_reg_16_23_inst : DFFR_X1 port map( D => n6837, CK => CLK, RN => 
                           n3209, Q => REGISTERS_16_23_port, QN => n_2124);
   REGISTERS_reg_16_22_inst : DFFR_X1 port map( D => n6838, CK => CLK, RN => 
                           n3209, Q => REGISTERS_16_22_port, QN => n_2125);
   REGISTERS_reg_16_21_inst : DFFR_X1 port map( D => n6839, CK => CLK, RN => 
                           n3209, Q => REGISTERS_16_21_port, QN => n_2126);
   REGISTERS_reg_16_20_inst : DFFR_X1 port map( D => n6840, CK => CLK, RN => 
                           n3209, Q => REGISTERS_16_20_port, QN => n_2127);
   REGISTERS_reg_16_19_inst : DFFR_X1 port map( D => n6841, CK => CLK, RN => 
                           n3209, Q => REGISTERS_16_19_port, QN => n_2128);
   REGISTERS_reg_16_18_inst : DFFR_X1 port map( D => n6842, CK => CLK, RN => 
                           n3209, Q => REGISTERS_16_18_port, QN => n_2129);
   REGISTERS_reg_16_17_inst : DFFR_X1 port map( D => n6843, CK => CLK, RN => 
                           n3209, Q => REGISTERS_16_17_port, QN => n_2130);
   REGISTERS_reg_16_16_inst : DFFR_X1 port map( D => n6844, CK => CLK, RN => 
                           n3209, Q => REGISTERS_16_16_port, QN => n_2131);
   REGISTERS_reg_16_15_inst : DFFR_X1 port map( D => n6845, CK => CLK, RN => 
                           n3209, Q => REGISTERS_16_15_port, QN => n_2132);
   REGISTERS_reg_16_14_inst : DFFR_X1 port map( D => n6846, CK => CLK, RN => 
                           n3209, Q => REGISTERS_16_14_port, QN => n_2133);
   REGISTERS_reg_16_13_inst : DFFR_X1 port map( D => n6847, CK => CLK, RN => 
                           n3209, Q => REGISTERS_16_13_port, QN => n_2134);
   REGISTERS_reg_16_12_inst : DFFR_X1 port map( D => n6848, CK => CLK, RN => 
                           n3209, Q => REGISTERS_16_12_port, QN => n_2135);
   REGISTERS_reg_16_11_inst : DFFR_X1 port map( D => n6849, CK => CLK, RN => 
                           n3208, Q => REGISTERS_16_11_port, QN => n_2136);
   REGISTERS_reg_16_10_inst : DFFR_X1 port map( D => n6850, CK => CLK, RN => 
                           n3208, Q => REGISTERS_16_10_port, QN => n_2137);
   REGISTERS_reg_16_9_inst : DFFR_X1 port map( D => n6851, CK => CLK, RN => 
                           n3208, Q => REGISTERS_16_9_port, QN => n_2138);
   REGISTERS_reg_16_8_inst : DFFR_X1 port map( D => n6852, CK => CLK, RN => 
                           n3208, Q => REGISTERS_16_8_port, QN => n_2139);
   REGISTERS_reg_16_7_inst : DFFR_X1 port map( D => n6853, CK => CLK, RN => 
                           n3208, Q => REGISTERS_16_7_port, QN => n_2140);
   REGISTERS_reg_16_6_inst : DFFR_X1 port map( D => n6854, CK => CLK, RN => 
                           n3208, Q => REGISTERS_16_6_port, QN => n_2141);
   REGISTERS_reg_16_5_inst : DFFR_X1 port map( D => n6855, CK => CLK, RN => 
                           n3208, Q => REGISTERS_16_5_port, QN => n_2142);
   REGISTERS_reg_16_4_inst : DFFR_X1 port map( D => n6856, CK => CLK, RN => 
                           n3208, Q => REGISTERS_16_4_port, QN => n_2143);
   REGISTERS_reg_16_3_inst : DFFR_X1 port map( D => n6857, CK => CLK, RN => 
                           n3208, Q => REGISTERS_16_3_port, QN => n_2144);
   REGISTERS_reg_16_2_inst : DFFR_X1 port map( D => n6858, CK => CLK, RN => 
                           n3208, Q => REGISTERS_16_2_port, QN => n_2145);
   REGISTERS_reg_16_1_inst : DFFR_X1 port map( D => n6859, CK => CLK, RN => 
                           n3208, Q => REGISTERS_16_1_port, QN => n_2146);
   REGISTERS_reg_16_0_inst : DFFR_X1 port map( D => n6860, CK => CLK, RN => 
                           n3208, Q => REGISTERS_16_0_port, QN => n_2147);
   REGISTERS_reg_12_31_inst : DFFR_X1 port map( D => n6701, CK => CLK, RN => 
                           n3225, Q => REGISTERS_12_31_port, QN => n_2148);
   REGISTERS_reg_12_30_inst : DFFR_X1 port map( D => n6702, CK => CLK, RN => 
                           n3225, Q => REGISTERS_12_30_port, QN => n_2149);
   REGISTERS_reg_12_29_inst : DFFR_X1 port map( D => n6703, CK => CLK, RN => 
                           n3225, Q => REGISTERS_12_29_port, QN => n_2150);
   REGISTERS_reg_12_28_inst : DFFR_X1 port map( D => n6704, CK => CLK, RN => 
                           n3225, Q => REGISTERS_12_28_port, QN => n_2151);
   REGISTERS_reg_12_27_inst : DFFR_X1 port map( D => n6705, CK => CLK, RN => 
                           n3224, Q => REGISTERS_12_27_port, QN => n_2152);
   REGISTERS_reg_12_26_inst : DFFR_X1 port map( D => n6706, CK => CLK, RN => 
                           n3224, Q => REGISTERS_12_26_port, QN => n_2153);
   REGISTERS_reg_12_25_inst : DFFR_X1 port map( D => n6707, CK => CLK, RN => 
                           n3224, Q => REGISTERS_12_25_port, QN => n_2154);
   REGISTERS_reg_12_24_inst : DFFR_X1 port map( D => n6708, CK => CLK, RN => 
                           n3224, Q => REGISTERS_12_24_port, QN => n_2155);
   REGISTERS_reg_12_23_inst : DFFR_X1 port map( D => n6709, CK => CLK, RN => 
                           n3224, Q => REGISTERS_12_23_port, QN => n_2156);
   REGISTERS_reg_12_22_inst : DFFR_X1 port map( D => n6710, CK => CLK, RN => 
                           n3224, Q => REGISTERS_12_22_port, QN => n_2157);
   REGISTERS_reg_12_21_inst : DFFR_X1 port map( D => n6711, CK => CLK, RN => 
                           n3224, Q => REGISTERS_12_21_port, QN => n_2158);
   REGISTERS_reg_12_20_inst : DFFR_X1 port map( D => n6712, CK => CLK, RN => 
                           n3224, Q => REGISTERS_12_20_port, QN => n_2159);
   REGISTERS_reg_12_19_inst : DFFR_X1 port map( D => n6713, CK => CLK, RN => 
                           n3224, Q => REGISTERS_12_19_port, QN => n_2160);
   REGISTERS_reg_12_18_inst : DFFR_X1 port map( D => n6714, CK => CLK, RN => 
                           n3224, Q => REGISTERS_12_18_port, QN => n_2161);
   REGISTERS_reg_12_17_inst : DFFR_X1 port map( D => n6715, CK => CLK, RN => 
                           n3224, Q => REGISTERS_12_17_port, QN => n_2162);
   REGISTERS_reg_12_16_inst : DFFR_X1 port map( D => n6716, CK => CLK, RN => 
                           n3224, Q => REGISTERS_12_16_port, QN => n_2163);
   REGISTERS_reg_12_15_inst : DFFR_X1 port map( D => n6717, CK => CLK, RN => 
                           n3223, Q => REGISTERS_12_15_port, QN => n_2164);
   REGISTERS_reg_12_14_inst : DFFR_X1 port map( D => n6718, CK => CLK, RN => 
                           n3223, Q => REGISTERS_12_14_port, QN => n_2165);
   REGISTERS_reg_12_13_inst : DFFR_X1 port map( D => n6719, CK => CLK, RN => 
                           n3223, Q => REGISTERS_12_13_port, QN => n_2166);
   REGISTERS_reg_12_12_inst : DFFR_X1 port map( D => n6720, CK => CLK, RN => 
                           n3223, Q => REGISTERS_12_12_port, QN => n_2167);
   REGISTERS_reg_12_11_inst : DFFR_X1 port map( D => n6721, CK => CLK, RN => 
                           n3223, Q => REGISTERS_12_11_port, QN => n_2168);
   REGISTERS_reg_12_10_inst : DFFR_X1 port map( D => n6722, CK => CLK, RN => 
                           n3223, Q => REGISTERS_12_10_port, QN => n_2169);
   REGISTERS_reg_12_9_inst : DFFR_X1 port map( D => n6723, CK => CLK, RN => 
                           n3223, Q => REGISTERS_12_9_port, QN => n_2170);
   REGISTERS_reg_12_8_inst : DFFR_X1 port map( D => n6724, CK => CLK, RN => 
                           n3223, Q => REGISTERS_12_8_port, QN => n_2171);
   REGISTERS_reg_12_7_inst : DFFR_X1 port map( D => n6725, CK => CLK, RN => 
                           n3223, Q => REGISTERS_12_7_port, QN => n_2172);
   REGISTERS_reg_12_6_inst : DFFR_X1 port map( D => n6726, CK => CLK, RN => 
                           n3223, Q => REGISTERS_12_6_port, QN => n_2173);
   REGISTERS_reg_12_5_inst : DFFR_X1 port map( D => n6727, CK => CLK, RN => 
                           n3223, Q => REGISTERS_12_5_port, QN => n_2174);
   REGISTERS_reg_12_4_inst : DFFR_X1 port map( D => n6728, CK => CLK, RN => 
                           n3223, Q => REGISTERS_12_4_port, QN => n_2175);
   REGISTERS_reg_12_3_inst : DFFR_X1 port map( D => n6729, CK => CLK, RN => 
                           n3221, Q => REGISTERS_12_3_port, QN => n_2176);
   REGISTERS_reg_12_2_inst : DFFR_X1 port map( D => n6730, CK => CLK, RN => 
                           n3221, Q => REGISTERS_12_2_port, QN => n_2177);
   REGISTERS_reg_12_1_inst : DFFR_X1 port map( D => n6731, CK => CLK, RN => 
                           n3221, Q => REGISTERS_12_1_port, QN => n_2178);
   REGISTERS_reg_12_0_inst : DFFR_X1 port map( D => n6732, CK => CLK, RN => 
                           n3221, Q => REGISTERS_12_0_port, QN => n_2179);
   REGISTERS_reg_11_31_inst : DFFR_X1 port map( D => n6669, CK => CLK, RN => 
                           n3228, Q => REGISTERS_11_31_port, QN => n_2180);
   REGISTERS_reg_11_30_inst : DFFR_X1 port map( D => n6670, CK => CLK, RN => 
                           n3228, Q => REGISTERS_11_30_port, QN => n_2181);
   REGISTERS_reg_11_29_inst : DFFR_X1 port map( D => n6671, CK => CLK, RN => 
                           n3228, Q => REGISTERS_11_29_port, QN => n_2182);
   REGISTERS_reg_11_28_inst : DFFR_X1 port map( D => n6672, CK => CLK, RN => 
                           n3228, Q => REGISTERS_11_28_port, QN => n_2183);
   REGISTERS_reg_11_27_inst : DFFR_X1 port map( D => n6673, CK => CLK, RN => 
                           n3228, Q => REGISTERS_11_27_port, QN => n_2184);
   REGISTERS_reg_11_26_inst : DFFR_X1 port map( D => n6674, CK => CLK, RN => 
                           n3228, Q => REGISTERS_11_26_port, QN => n_2185);
   REGISTERS_reg_11_25_inst : DFFR_X1 port map( D => n6675, CK => CLK, RN => 
                           n3228, Q => REGISTERS_11_25_port, QN => n_2186);
   REGISTERS_reg_11_24_inst : DFFR_X1 port map( D => n6676, CK => CLK, RN => 
                           n3228, Q => REGISTERS_11_24_port, QN => n_2187);
   REGISTERS_reg_11_23_inst : DFFR_X1 port map( D => n6677, CK => CLK, RN => 
                           n3228, Q => REGISTERS_11_23_port, QN => n_2188);
   REGISTERS_reg_11_22_inst : DFFR_X1 port map( D => n6678, CK => CLK, RN => 
                           n3228, Q => REGISTERS_11_22_port, QN => n_2189);
   REGISTERS_reg_11_21_inst : DFFR_X1 port map( D => n6679, CK => CLK, RN => 
                           n3228, Q => REGISTERS_11_21_port, QN => n_2190);
   REGISTERS_reg_11_20_inst : DFFR_X1 port map( D => n6680, CK => CLK, RN => 
                           n3228, Q => REGISTERS_11_20_port, QN => n_2191);
   REGISTERS_reg_11_19_inst : DFFR_X1 port map( D => n6681, CK => CLK, RN => 
                           n3227, Q => REGISTERS_11_19_port, QN => n_2192);
   REGISTERS_reg_11_18_inst : DFFR_X1 port map( D => n6682, CK => CLK, RN => 
                           n3227, Q => REGISTERS_11_18_port, QN => n_2193);
   REGISTERS_reg_11_17_inst : DFFR_X1 port map( D => n6683, CK => CLK, RN => 
                           n3227, Q => REGISTERS_11_17_port, QN => n_2194);
   REGISTERS_reg_11_16_inst : DFFR_X1 port map( D => n6684, CK => CLK, RN => 
                           n3227, Q => REGISTERS_11_16_port, QN => n_2195);
   REGISTERS_reg_11_15_inst : DFFR_X1 port map( D => n6685, CK => CLK, RN => 
                           n3227, Q => REGISTERS_11_15_port, QN => n_2196);
   REGISTERS_reg_11_14_inst : DFFR_X1 port map( D => n6686, CK => CLK, RN => 
                           n3227, Q => REGISTERS_11_14_port, QN => n_2197);
   REGISTERS_reg_11_13_inst : DFFR_X1 port map( D => n6687, CK => CLK, RN => 
                           n3227, Q => REGISTERS_11_13_port, QN => n_2198);
   REGISTERS_reg_11_12_inst : DFFR_X1 port map( D => n6688, CK => CLK, RN => 
                           n3227, Q => REGISTERS_11_12_port, QN => n_2199);
   REGISTERS_reg_11_11_inst : DFFR_X1 port map( D => n6689, CK => CLK, RN => 
                           n3227, Q => REGISTERS_11_11_port, QN => n_2200);
   REGISTERS_reg_11_10_inst : DFFR_X1 port map( D => n6690, CK => CLK, RN => 
                           n3227, Q => REGISTERS_11_10_port, QN => n_2201);
   REGISTERS_reg_11_9_inst : DFFR_X1 port map( D => n6691, CK => CLK, RN => 
                           n3227, Q => REGISTERS_11_9_port, QN => n_2202);
   REGISTERS_reg_11_8_inst : DFFR_X1 port map( D => n6692, CK => CLK, RN => 
                           n3227, Q => REGISTERS_11_8_port, QN => n_2203);
   REGISTERS_reg_11_7_inst : DFFR_X1 port map( D => n6693, CK => CLK, RN => 
                           n3225, Q => REGISTERS_11_7_port, QN => n_2204);
   REGISTERS_reg_11_6_inst : DFFR_X1 port map( D => n6694, CK => CLK, RN => 
                           n3225, Q => REGISTERS_11_6_port, QN => n_2205);
   REGISTERS_reg_11_5_inst : DFFR_X1 port map( D => n6695, CK => CLK, RN => 
                           n3225, Q => REGISTERS_11_5_port, QN => n_2206);
   REGISTERS_reg_11_4_inst : DFFR_X1 port map( D => n6696, CK => CLK, RN => 
                           n3225, Q => REGISTERS_11_4_port, QN => n_2207);
   REGISTERS_reg_11_3_inst : DFFR_X1 port map( D => n6697, CK => CLK, RN => 
                           n3225, Q => REGISTERS_11_3_port, QN => n_2208);
   REGISTERS_reg_11_2_inst : DFFR_X1 port map( D => n6698, CK => CLK, RN => 
                           n3225, Q => REGISTERS_11_2_port, QN => n_2209);
   REGISTERS_reg_11_1_inst : DFFR_X1 port map( D => n6699, CK => CLK, RN => 
                           n3225, Q => REGISTERS_11_1_port, QN => n_2210);
   REGISTERS_reg_11_0_inst : DFFR_X1 port map( D => n6700, CK => CLK, RN => 
                           n3225, Q => REGISTERS_11_0_port, QN => n_2211);
   CWP_reg_6_inst : DFFR_X1 port map( D => n9133, CK => CLK, RN => n2970, Q => 
                           CWP_6_port, QN => n2898);
   CWP_reg_5_inst : DFFR_X1 port map( D => n9134, CK => CLK, RN => n2969, Q => 
                           CWP_5_port, QN => n2916);
   CWP_reg_4_inst : DFFR_X1 port map( D => n9135, CK => CLK, RN => n2968, Q => 
                           CWP_4_port, QN => N8791);
   CWP_reg_3_inst : DFFR_X1 port map( D => n9136, CK => CLK, RN => n2967, Q => 
                           N8790, QN => n2918);
   CWP_reg_2_inst : DFFR_X1 port map( D => n9137, CK => CLK, RN => n2966, Q => 
                           N8789, QN => n2919);
   CWP_reg_1_inst : DFFR_X1 port map( D => n9138, CK => CLK, RN => n2965, Q => 
                           N8788, QN => n2920);
   CWP_reg_0_inst : DFFR_X1 port map( D => n9139, CK => CLK, RN => n2964, Q => 
                           N8787, QN => n2921);
   U3 : AOI22_X1 port map( A1 => N8430, A2 => n10918, B1 => N8423, B2 => N8415,
                           ZN => n6266);
   U4 : AOI22_X1 port map( A1 => N8574, A2 => n10919, B1 => N8567, B2 => N8559,
                           ZN => n4823);
   U5 : NOR2_X1 port map( A1 => n3378, A2 => n6314, ZN => n6249);
   U6 : NOR2_X1 port map( A1 => n3387, A2 => n4871, ZN => n4806);
   U7 : AOI22_X1 port map( A1 => N2165, A2 => n3391, B1 => N2158, B2 => N2151, 
                           ZN => n3108);
   U8 : AOI22_X1 port map( A1 => N2166, A2 => n3391, B1 => N2159, B2 => N2151, 
                           ZN => n3107);
   U9 : XOR2_X1 port map( A => CWP_5_port, B => CWP_4_port, Z => n1);
   U10 : NOR2_X1 port map( A1 => n3378, A2 => n3379, ZN => n6247);
   U11 : NOR2_X1 port map( A1 => n3387, A2 => n3388, ZN => n4804);
   U12 : NAND4_X1 port map( A1 => n3106, A2 => n3107, A3 => n3108, A4 => n3109,
                           ZN => n3029);
   U13 : NAND4_X1 port map( A1 => n3106, A2 => n3108, A3 => n3109, A4 => n3365,
                           ZN => n3309);
   U14 : NAND4_X1 port map( A1 => n3106, A2 => n3107, A3 => n3109, A4 => n3366,
                           ZN => n3179);
   U15 : NAND4_X1 port map( A1 => n3106, A2 => n3107, A3 => n3368, A4 => n3366,
                           ZN => n3244);
   U16 : NAND4_X1 port map( A1 => n3106, A2 => n3107, A3 => n3108, A4 => n3368,
                           ZN => n3114);
   U17 : NOR2_X1 port map( A1 => n6265, A2 => n6264, ZN => n6296);
   U18 : NOR2_X1 port map( A1 => n4822, A2 => n4821, ZN => n4853);
   U20 : NOR2_X1 port map( A1 => n3376, A2 => n6264, ZN => n6283);
   U21 : NOR2_X1 port map( A1 => n3385, A2 => n4821, ZN => n4840);
   U22 : NOR2_X1 port map( A1 => n6314, A2 => n6315, ZN => n6251);
   U24 : NOR2_X1 port map( A1 => n4871, A2 => n4872, ZN => n4808);
   U25 : NOR2_X1 port map( A1 => n3379, A2 => n6315, ZN => n6250);
   U26 : NOR2_X1 port map( A1 => n3388, A2 => n4872, ZN => n4807);
   U27 : INV_X1 port map( A => N2166, ZN => N2165);
   U28 : BUF_X1 port map( A => n3345, Z => n3301);
   U30 : BUF_X1 port map( A => n3347, Z => n3300);
   U31 : BUF_X1 port map( A => n3347, Z => n3298);
   U32 : BUF_X1 port map( A => n3347, Z => n3297);
   U33 : BUF_X1 port map( A => n3349, Z => n3296);
   U34 : BUF_X1 port map( A => n3349, Z => n3293);
   U35 : BUF_X1 port map( A => n3350, Z => n3292);
   U36 : BUF_X1 port map( A => n3350, Z => n3290);
   U37 : BUF_X1 port map( A => n3350, Z => n3289);
   U38 : BUF_X1 port map( A => n3352, Z => n3288);
   U39 : BUF_X1 port map( A => n3349, Z => n3294);
   U40 : BUF_X1 port map( A => n3334, Z => n3331);
   U41 : BUF_X1 port map( A => n3334, Z => n3330);
   U42 : BUF_X1 port map( A => n3335, Z => n3329);
   U43 : BUF_X1 port map( A => n3335, Z => n3327);
   U44 : BUF_X1 port map( A => n3335, Z => n3326);
   U45 : BUF_X1 port map( A => n3337, Z => n3325);
   U46 : BUF_X1 port map( A => n3337, Z => n3323);
   U47 : BUF_X1 port map( A => n3337, Z => n3322);
   U48 : BUF_X1 port map( A => n3338, Z => n3321);
   U49 : BUF_X1 port map( A => n3338, Z => n3319);
   U50 : BUF_X1 port map( A => n3339, Z => n3317);
   U51 : BUF_X1 port map( A => n3339, Z => n3315);
   U52 : BUF_X1 port map( A => n3339, Z => n3314);
   U53 : BUF_X1 port map( A => n3341, Z => n3313);
   U54 : BUF_X1 port map( A => n3341, Z => n3311);
   U55 : BUF_X1 port map( A => n3341, Z => n3310);
   U56 : BUF_X1 port map( A => n3344, Z => n3308);
   U57 : BUF_X1 port map( A => n3344, Z => n3306);
   U58 : BUF_X1 port map( A => n3344, Z => n3305);
   U59 : BUF_X1 port map( A => n3345, Z => n3304);
   U60 : BUF_X1 port map( A => n3338, Z => n3318);
   U61 : BUF_X1 port map( A => n3352, Z => n3286);
   U62 : BUF_X1 port map( A => n3361, Z => n3265);
   U63 : BUF_X1 port map( A => n3355, Z => n3277);
   U64 : BUF_X1 port map( A => n3361, Z => n3266);
   U65 : BUF_X1 port map( A => n3355, Z => n3278);
   U66 : BUF_X1 port map( A => n3361, Z => n3268);
   U67 : BUF_X1 port map( A => n3355, Z => n3280);
   U68 : BUF_X1 port map( A => n3360, Z => n3269);
   U69 : BUF_X1 port map( A => n3354, Z => n3281);
   U70 : BUF_X1 port map( A => n3360, Z => n3270);
   U71 : BUF_X1 port map( A => n3354, Z => n3282);
   U72 : BUF_X1 port map( A => n3360, Z => n3272);
   U73 : BUF_X1 port map( A => n3354, Z => n3284);
   U74 : BUF_X1 port map( A => n3357, Z => n3273);
   U75 : BUF_X1 port map( A => n3352, Z => n3285);
   U76 : BUF_X1 port map( A => n3357, Z => n3274);
   U77 : BUF_X1 port map( A => n3357, Z => n3276);
   U78 : BUF_X1 port map( A => n3345, Z => n3302);
   U79 : BUF_X1 port map( A => n3334, Z => n3333);
   U80 : BUF_X1 port map( A => n4887, Z => n716);
   U81 : BUF_X1 port map( A => n3444, Z => n1428);
   U82 : BUF_X1 port map( A => n4887, Z => n717);
   U83 : BUF_X1 port map( A => n3444, Z => n1429);
   U84 : BUF_X1 port map( A => n4888, Z => n713);
   U85 : BUF_X1 port map( A => n3445, Z => n1425);
   U86 : BUF_X1 port map( A => n4888, Z => n714);
   U87 : BUF_X1 port map( A => n3445, Z => n1426);
   U88 : BUF_X1 port map( A => n4887, Z => n718);
   U89 : BUF_X1 port map( A => n3444, Z => n1430);
   U90 : BUF_X1 port map( A => n4957, Z => n464);
   U91 : BUF_X1 port map( A => n3514, Z => n1176);
   U92 : BUF_X1 port map( A => n4957, Z => n465);
   U93 : BUF_X1 port map( A => n3514, Z => n1177);
   U94 : BUF_X1 port map( A => n4927, Z => n623);
   U95 : BUF_X1 port map( A => n4964, Z => n446);
   U96 : BUF_X1 port map( A => n4995, Z => n28);
   U97 : BUF_X1 port map( A => n3484, Z => n1335);
   U98 : BUF_X1 port map( A => n3521, Z => n1158);
   U99 : BUF_X1 port map( A => n3552, Z => n740);
   U100 : BUF_X1 port map( A => n4927, Z => n624);
   U101 : BUF_X1 port map( A => n4964, Z => n447);
   U102 : BUF_X1 port map( A => n4995, Z => n29);
   U103 : BUF_X1 port map( A => n3484, Z => n1336);
   U104 : BUF_X1 port map( A => n3521, Z => n1159);
   U105 : BUF_X1 port map( A => n3552, Z => n741);
   U106 : BUF_X1 port map( A => n4888, Z => n715);
   U107 : BUF_X1 port map( A => n3445, Z => n1427);
   U108 : BUF_X1 port map( A => n4909, Z => n654);
   U109 : BUF_X1 port map( A => n3466, Z => n1366);
   U110 : BUF_X1 port map( A => n4909, Z => n653);
   U111 : BUF_X1 port map( A => n3466, Z => n1365);
   U112 : BUF_X1 port map( A => n4957, Z => n466);
   U113 : BUF_X1 port map( A => n3514, Z => n1178);
   U114 : BUF_X1 port map( A => n4927, Z => n625);
   U115 : BUF_X1 port map( A => n4964, Z => n448);
   U116 : BUF_X1 port map( A => n4995, Z => n30);
   U117 : BUF_X1 port map( A => n3484, Z => n1337);
   U118 : BUF_X1 port map( A => n3521, Z => n1160);
   U119 : BUF_X1 port map( A => n3552, Z => n742);
   U120 : BUF_X1 port map( A => n4909, Z => n655);
   U121 : BUF_X1 port map( A => n3466, Z => n1367);
   U122 : BUF_X1 port map( A => n3354, Z => n3361);
   U123 : BUF_X1 port map( A => n3363, Z => n3355);
   U124 : BUF_X1 port map( A => n3352, Z => n3360);
   U125 : BUF_X1 port map( A => n3347, Z => n3354);
   U126 : BUF_X1 port map( A => n3349, Z => n3357);
   U127 : BUF_X1 port map( A => n3363, Z => n3347);
   U128 : BUF_X1 port map( A => n3363, Z => n3350);
   U129 : BUF_X1 port map( A => n3363, Z => n3349);
   U130 : BUF_X1 port map( A => n3341, Z => n3337);
   U131 : BUF_X1 port map( A => n3344, Z => n3339);
   U132 : BUF_X1 port map( A => n3333, Z => n3341);
   U133 : BUF_X1 port map( A => n3333, Z => n3344);
   U134 : BUF_X1 port map( A => n3335, Z => n3338);
   U135 : BUF_X1 port map( A => n3350, Z => n3352);
   U136 : BUF_X1 port map( A => n3334, Z => n3345);
   U137 : BUF_X1 port map( A => n3355, Z => n3334);
   U138 : BUF_X1 port map( A => n3361, Z => n3335);
   U139 : NAND2_X1 port map( A1 => n3383, A2 => n3343, ZN => n3030);
   U140 : BUF_X1 port map( A => n4980, Z => n70);
   U141 : BUF_X1 port map( A => n3537, Z => n782);
   U142 : BUF_X1 port map( A => n4980, Z => n71);
   U143 : BUF_X1 port map( A => n3537, Z => n783);
   U144 : BUF_X1 port map( A => n4918, Z => n650);
   U145 : BUF_X1 port map( A => n3475, Z => n1362);
   U146 : BUF_X1 port map( A => n4918, Z => n651);
   U147 : BUF_X1 port map( A => n3475, Z => n1363);
   U148 : BUF_X1 port map( A => n4949, Z => n488);
   U149 : BUF_X1 port map( A => n3506, Z => n1296);
   U150 : BUF_X1 port map( A => n4949, Z => n489);
   U151 : BUF_X1 port map( A => n3506, Z => n1297);
   U152 : BUF_X1 port map( A => n4919, Z => n647);
   U153 : BUF_X1 port map( A => n3476, Z => n1359);
   U154 : BUF_X1 port map( A => n4919, Z => n648);
   U155 : BUF_X1 port map( A => n3476, Z => n1360);
   U156 : BUF_X1 port map( A => n4950, Z => n485);
   U157 : BUF_X1 port map( A => n4981, Z => n67);
   U158 : BUF_X1 port map( A => n3507, Z => n1197);
   U159 : BUF_X1 port map( A => n3538, Z => n779);
   U160 : BUF_X1 port map( A => n4950, Z => n486);
   U161 : BUF_X1 port map( A => n4981, Z => n68);
   U162 : BUF_X1 port map( A => n3507, Z => n1198);
   U163 : BUF_X1 port map( A => n3538, Z => n780);
   U164 : BUF_X1 port map( A => n4898, Z => n683);
   U165 : BUF_X1 port map( A => n4929, Z => n617);
   U166 : BUF_X1 port map( A => n4960, Z => n455);
   U167 : BUF_X1 port map( A => n4991, Z => n37);
   U168 : BUF_X1 port map( A => n3455, Z => n1395);
   U169 : BUF_X1 port map( A => n3486, Z => n1329);
   U170 : BUF_X1 port map( A => n3517, Z => n1167);
   U171 : BUF_X1 port map( A => n3548, Z => n749);
   U172 : BUF_X1 port map( A => n4898, Z => n684);
   U173 : BUF_X1 port map( A => n4929, Z => n618);
   U174 : BUF_X1 port map( A => n4960, Z => n456);
   U175 : BUF_X1 port map( A => n4991, Z => n38);
   U176 : BUF_X1 port map( A => n3455, Z => n1396);
   U177 : BUF_X1 port map( A => n3486, Z => n1330);
   U178 : BUF_X1 port map( A => n3517, Z => n1168);
   U179 : BUF_X1 port map( A => n3548, Z => n750);
   U180 : BUF_X1 port map( A => n4904, Z => n668);
   U181 : BUF_X1 port map( A => n4907, Z => n659);
   U182 : BUF_X1 port map( A => n4935, Z => n602);
   U183 : BUF_X1 port map( A => n4938, Z => n593);
   U184 : BUF_X1 port map( A => n4966, Z => n440);
   U185 : BUF_X1 port map( A => n4969, Z => n79);
   U186 : BUF_X1 port map( A => n4997, Z => n22);
   U187 : BUF_X1 port map( A => n5000, Z => n12);
   U188 : BUF_X1 port map( A => n3461, Z => n1380);
   U189 : BUF_X1 port map( A => n3464, Z => n1371);
   U190 : BUF_X1 port map( A => n3492, Z => n1314);
   U191 : BUF_X1 port map( A => n3495, Z => n1305);
   U192 : BUF_X1 port map( A => n3523, Z => n1152);
   U194 : BUF_X1 port map( A => n3526, Z => n1143);
   U195 : BUF_X1 port map( A => n3554, Z => n734);
   U196 : BUF_X1 port map( A => n3557, Z => n725);
   U197 : BUF_X1 port map( A => n4904, Z => n669);
   U198 : BUF_X1 port map( A => n4907, Z => n660);
   U199 : BUF_X1 port map( A => n4935, Z => n603);
   U200 : BUF_X1 port map( A => n4938, Z => n594);
   U201 : BUF_X1 port map( A => n4966, Z => n441);
   U202 : BUF_X1 port map( A => n4969, Z => n432);
   U203 : BUF_X1 port map( A => n4997, Z => n23);
   U204 : BUF_X1 port map( A => n5000, Z => n13);
   U205 : BUF_X1 port map( A => n3461, Z => n1381);
   U206 : BUF_X1 port map( A => n3464, Z => n1372);
   U207 : BUF_X1 port map( A => n3492, Z => n1315);
   U208 : BUF_X1 port map( A => n3495, Z => n1306);
   U209 : BUF_X1 port map( A => n3523, Z => n1153);
   U210 : BUF_X1 port map( A => n3526, Z => n1144);
   U211 : BUF_X1 port map( A => n3554, Z => n735);
   U212 : BUF_X1 port map( A => n3557, Z => n726);
   U213 : BUF_X1 port map( A => n4899, Z => n680);
   U214 : BUF_X1 port map( A => n4930, Z => n614);
   U215 : BUF_X1 port map( A => n4961, Z => n452);
   U216 : BUF_X1 port map( A => n4992, Z => n34);
   U217 : BUF_X1 port map( A => n3456, Z => n1392);
   U218 : BUF_X1 port map( A => n3487, Z => n1326);
   U219 : BUF_X1 port map( A => n3518, Z => n1164);
   U220 : BUF_X1 port map( A => n3549, Z => n746);
   U221 : BUF_X1 port map( A => n4899, Z => n681);
   U222 : BUF_X1 port map( A => n4930, Z => n615);
   U223 : BUF_X1 port map( A => n4961, Z => n453);
   U224 : BUF_X1 port map( A => n4992, Z => n35);
   U225 : BUF_X1 port map( A => n3456, Z => n1393);
   U226 : BUF_X1 port map( A => n3487, Z => n1327);
   U228 : BUF_X1 port map( A => n3518, Z => n1165);
   U229 : BUF_X1 port map( A => n3549, Z => n747);
   U230 : BUF_X1 port map( A => n4891, Z => n704);
   U231 : BUF_X1 port map( A => n3448, Z => n1416);
   U232 : BUF_X1 port map( A => n4891, Z => n705);
   U233 : BUF_X1 port map( A => n3448, Z => n1417);
   U234 : BUF_X1 port map( A => n4990, Z => n40);
   U235 : BUF_X1 port map( A => n4996, Z => n25);
   U236 : BUF_X1 port map( A => n3547, Z => n752);
   U237 : BUF_X1 port map( A => n3553, Z => n737);
   U238 : BUF_X1 port map( A => n4990, Z => n41);
   U239 : BUF_X1 port map( A => n4996, Z => n26);
   U240 : BUF_X1 port map( A => n3547, Z => n753);
   U241 : BUF_X1 port map( A => n3553, Z => n738);
   U242 : BUF_X1 port map( A => n4894, Z => n695);
   U243 : BUF_X1 port map( A => n4897, Z => n686);
   U244 : BUF_X1 port map( A => n4903, Z => n671);
   U245 : BUF_X1 port map( A => n4922, Z => n638);
   U246 : BUF_X1 port map( A => n4925, Z => n629);
   U247 : BUF_X1 port map( A => n4928, Z => n620);
   U248 : BUF_X1 port map( A => n4934, Z => n605);
   U249 : BUF_X1 port map( A => n4953, Z => n476);
   U250 : BUF_X1 port map( A => n4956, Z => n467);
   U251 : BUF_X1 port map( A => n4959, Z => n458);
   U252 : BUF_X1 port map( A => n4965, Z => n443);
   U253 : BUF_X1 port map( A => n4984, Z => n58);
   U254 : BUF_X1 port map( A => n4987, Z => n49);
   U255 : BUF_X1 port map( A => n3451, Z => n1407);
   U256 : BUF_X1 port map( A => n3454, Z => n1398);
   U257 : BUF_X1 port map( A => n3460, Z => n1383);
   U258 : BUF_X1 port map( A => n3479, Z => n1350);
   U259 : BUF_X1 port map( A => n3482, Z => n1341);
   U260 : BUF_X1 port map( A => n3485, Z => n1332);
   U261 : BUF_X1 port map( A => n3491, Z => n1317);
   U262 : BUF_X1 port map( A => n3510, Z => n1188);
   U263 : BUF_X1 port map( A => n3513, Z => n1179);
   U264 : BUF_X1 port map( A => n3516, Z => n1170);
   U265 : BUF_X1 port map( A => n3522, Z => n1155);
   U266 : BUF_X1 port map( A => n3541, Z => n770);
   U267 : BUF_X1 port map( A => n3544, Z => n761);
   U268 : BUF_X1 port map( A => n4894, Z => n696);
   U269 : BUF_X1 port map( A => n4897, Z => n687);
   U270 : BUF_X1 port map( A => n4903, Z => n672);
   U271 : BUF_X1 port map( A => n4922, Z => n639);
   U272 : BUF_X1 port map( A => n4925, Z => n630);
   U273 : BUF_X1 port map( A => n4928, Z => n621);
   U274 : BUF_X1 port map( A => n4934, Z => n606);
   U275 : BUF_X1 port map( A => n4953, Z => n477);
   U276 : BUF_X1 port map( A => n4956, Z => n468);
   U277 : BUF_X1 port map( A => n4959, Z => n459);
   U278 : BUF_X1 port map( A => n4965, Z => n444);
   U279 : BUF_X1 port map( A => n4984, Z => n59);
   U280 : BUF_X1 port map( A => n4987, Z => n50);
   U281 : BUF_X1 port map( A => n3451, Z => n1408);
   U282 : BUF_X1 port map( A => n3454, Z => n1399);
   U283 : BUF_X1 port map( A => n3460, Z => n1384);
   U284 : BUF_X1 port map( A => n3479, Z => n1351);
   U285 : BUF_X1 port map( A => n3482, Z => n1342);
   U286 : BUF_X1 port map( A => n3485, Z => n1333);
   U287 : BUF_X1 port map( A => n3491, Z => n1318);
   U288 : BUF_X1 port map( A => n3510, Z => n1189);
   U289 : BUF_X1 port map( A => n3513, Z => n1180);
   U290 : BUF_X1 port map( A => n3516, Z => n1171);
   U291 : BUF_X1 port map( A => n3522, Z => n1156);
   U292 : BUF_X1 port map( A => n3541, Z => n771);
   U293 : BUF_X1 port map( A => n3544, Z => n762);
   U294 : BUF_X1 port map( A => n4980, Z => n72);
   U295 : BUF_X1 port map( A => n3537, Z => n1136);
   U296 : BUF_X1 port map( A => n4918, Z => n652);
   U297 : BUF_X1 port map( A => n3475, Z => n1364);
   U298 : BUF_X1 port map( A => n4949, Z => n490);
   U299 : BUF_X1 port map( A => n3506, Z => n1298);
   U300 : BUF_X1 port map( A => n4905, Z => n666);
   U301 : BUF_X1 port map( A => n4908, Z => n657);
   U302 : BUF_X1 port map( A => n4936, Z => n600);
   U303 : BUF_X1 port map( A => n4939, Z => n495);
   U304 : BUF_X1 port map( A => n4967, Z => n438);
   U305 : BUF_X1 port map( A => n4970, Z => n77);
   U306 : BUF_X1 port map( A => n4998, Z => n20);
   U307 : BUF_X1 port map( A => n5001, Z => n9);
   U308 : BUF_X1 port map( A => n3462, Z => n1378);
   U309 : BUF_X1 port map( A => n3465, Z => n1369);
   U310 : BUF_X1 port map( A => n3493, Z => n1312);
   U311 : BUF_X1 port map( A => n3496, Z => n1303);
   U312 : BUF_X1 port map( A => n3524, Z => n1150);
   U313 : BUF_X1 port map( A => n3527, Z => n1141);
   U314 : BUF_X1 port map( A => n3555, Z => n732);
   U315 : BUF_X1 port map( A => n3558, Z => n723);
   U316 : BUF_X1 port map( A => n4905, Z => n665);
   U317 : BUF_X1 port map( A => n4908, Z => n656);
   U318 : BUF_X1 port map( A => n4936, Z => n599);
   U319 : BUF_X1 port map( A => n4939, Z => n494);
   U320 : BUF_X1 port map( A => n4967, Z => n437);
   U321 : BUF_X1 port map( A => n4970, Z => n76);
   U322 : BUF_X1 port map( A => n4998, Z => n19);
   U323 : BUF_X1 port map( A => n5001, Z => n8);
   U324 : BUF_X1 port map( A => n3462, Z => n1377);
   U325 : BUF_X1 port map( A => n3465, Z => n1368);
   U326 : BUF_X1 port map( A => n3493, Z => n1311);
   U327 : BUF_X1 port map( A => n3496, Z => n1302);
   U328 : BUF_X1 port map( A => n3524, Z => n1149);
   U329 : BUF_X1 port map( A => n3527, Z => n1140);
   U330 : BUF_X1 port map( A => n3555, Z => n731);
   U331 : BUF_X1 port map( A => n3558, Z => n722);
   U332 : BUF_X1 port map( A => n4889, Z => n710);
   U333 : BUF_X1 port map( A => n3446, Z => n1422);
   U334 : BUF_X1 port map( A => n4889, Z => n711);
   U335 : BUF_X1 port map( A => n3446, Z => n1423);
   U336 : BUF_X1 port map( A => n4985, Z => n55);
   U337 : BUF_X1 port map( A => n4988, Z => n46);
   U338 : BUF_X1 port map( A => n3542, Z => n767);
   U339 : BUF_X1 port map( A => n3545, Z => n758);
   U340 : BUF_X1 port map( A => n4985, Z => n56);
   U341 : BUF_X1 port map( A => n4988, Z => n47);
   U342 : BUF_X1 port map( A => n3542, Z => n768);
   U343 : BUF_X1 port map( A => n3545, Z => n759);
   U344 : BUF_X1 port map( A => n4892, Z => n701);
   U345 : BUF_X1 port map( A => n3449, Z => n1413);
   U346 : BUF_X1 port map( A => n4892, Z => n702);
   U347 : BUF_X1 port map( A => n3449, Z => n1414);
   U348 : BUF_X1 port map( A => n4895, Z => n692);
   U349 : BUF_X1 port map( A => n4901, Z => n677);
   U350 : BUF_X1 port map( A => n4920, Z => n644);
   U351 : BUF_X1 port map( A => n4923, Z => n635);
   U352 : BUF_X1 port map( A => n4926, Z => n626);
   U353 : BUF_X1 port map( A => n4932, Z => n611);
   U354 : BUF_X1 port map( A => n4951, Z => n482);
   U355 : BUF_X1 port map( A => n4954, Z => n473);
   U356 : BUF_X1 port map( A => n4963, Z => n449);
   U357 : BUF_X1 port map( A => n4982, Z => n64);
   U358 : BUF_X1 port map( A => n4994, Z => n31);
   U359 : BUF_X1 port map( A => n3452, Z => n1404);
   U360 : BUF_X1 port map( A => n3458, Z => n1389);
   U361 : BUF_X1 port map( A => n3477, Z => n1356);
   U362 : BUF_X1 port map( A => n3480, Z => n1347);
   U363 : BUF_X1 port map( A => n3483, Z => n1338);
   U364 : BUF_X1 port map( A => n3489, Z => n1323);
   U365 : BUF_X1 port map( A => n3508, Z => n1194);
   U366 : BUF_X1 port map( A => n3511, Z => n1185);
   U367 : BUF_X1 port map( A => n3520, Z => n1161);
   U368 : BUF_X1 port map( A => n3539, Z => n776);
   U369 : BUF_X1 port map( A => n3551, Z => n743);
   U370 : BUF_X1 port map( A => n4895, Z => n693);
   U371 : BUF_X1 port map( A => n4901, Z => n678);
   U372 : BUF_X1 port map( A => n4920, Z => n645);
   U373 : BUF_X1 port map( A => n4923, Z => n636);
   U374 : BUF_X1 port map( A => n4926, Z => n627);
   U375 : BUF_X1 port map( A => n4932, Z => n612);
   U376 : BUF_X1 port map( A => n4951, Z => n483);
   U377 : BUF_X1 port map( A => n4954, Z => n474);
   U378 : BUF_X1 port map( A => n4963, Z => n450);
   U379 : BUF_X1 port map( A => n4982, Z => n65);
   U380 : BUF_X1 port map( A => n4994, Z => n32);
   U381 : BUF_X1 port map( A => n3452, Z => n1405);
   U382 : BUF_X1 port map( A => n3458, Z => n1390);
   U383 : BUF_X1 port map( A => n3477, Z => n1357);
   U384 : BUF_X1 port map( A => n3480, Z => n1348);
   U385 : BUF_X1 port map( A => n3483, Z => n1339);
   U386 : BUF_X1 port map( A => n3489, Z => n1324);
   U387 : BUF_X1 port map( A => n3508, Z => n1195);
   U388 : BUF_X1 port map( A => n3511, Z => n1186);
   U389 : BUF_X1 port map( A => n3520, Z => n1162);
   U390 : BUF_X1 port map( A => n3539, Z => n777);
   U391 : BUF_X1 port map( A => n3551, Z => n744);
   U392 : BUF_X1 port map( A => n4986, Z => n52);
   U393 : BUF_X1 port map( A => n4989, Z => n43);
   U394 : BUF_X1 port map( A => n3543, Z => n764);
   U395 : BUF_X1 port map( A => n3546, Z => n755);
   U396 : BUF_X1 port map( A => n4986, Z => n53);
   U397 : BUF_X1 port map( A => n4989, Z => n44);
   U398 : BUF_X1 port map( A => n3543, Z => n765);
   U399 : BUF_X1 port map( A => n3546, Z => n756);
   U400 : BUF_X1 port map( A => n4890, Z => n707);
   U401 : BUF_X1 port map( A => n4893, Z => n698);
   U402 : BUF_X1 port map( A => n4983, Z => n61);
   U403 : BUF_X1 port map( A => n3540, Z => n773);
   U404 : BUF_X1 port map( A => n4893, Z => n699);
   U405 : BUF_X1 port map( A => n4983, Z => n62);
   U406 : BUF_X1 port map( A => n3540, Z => n774);
   U407 : BUF_X1 port map( A => n4896, Z => n689);
   U408 : BUF_X1 port map( A => n4902, Z => n674);
   U409 : BUF_X1 port map( A => n4921, Z => n641);
   U410 : BUF_X1 port map( A => n4924, Z => n632);
   U411 : BUF_X1 port map( A => n4933, Z => n608);
   U412 : BUF_X1 port map( A => n4952, Z => n479);
   U413 : BUF_X1 port map( A => n4955, Z => n470);
   U414 : BUF_X1 port map( A => n4958, Z => n461);
   U415 : BUF_X1 port map( A => n3447, Z => n1419);
   U416 : BUF_X1 port map( A => n3450, Z => n1410);
   U417 : BUF_X1 port map( A => n3453, Z => n1401);
   U418 : BUF_X1 port map( A => n3459, Z => n1386);
   U419 : BUF_X1 port map( A => n3478, Z => n1353);
   U420 : BUF_X1 port map( A => n3481, Z => n1344);
   U421 : BUF_X1 port map( A => n3490, Z => n1320);
   U422 : BUF_X1 port map( A => n3509, Z => n1191);
   U423 : BUF_X1 port map( A => n3512, Z => n1182);
   U424 : BUF_X1 port map( A => n3515, Z => n1173);
   U425 : BUF_X1 port map( A => n4890, Z => n708);
   U426 : BUF_X1 port map( A => n4896, Z => n690);
   U427 : BUF_X1 port map( A => n4902, Z => n675);
   U428 : BUF_X1 port map( A => n4921, Z => n642);
   U429 : BUF_X1 port map( A => n4924, Z => n633);
   U430 : BUF_X1 port map( A => n4933, Z => n609);
   U431 : BUF_X1 port map( A => n4952, Z => n480);
   U432 : BUF_X1 port map( A => n4955, Z => n471);
   U433 : BUF_X1 port map( A => n4958, Z => n462);
   U434 : BUF_X1 port map( A => n3447, Z => n1420);
   U435 : BUF_X1 port map( A => n3450, Z => n1411);
   U436 : BUF_X1 port map( A => n3453, Z => n1402);
   U437 : BUF_X1 port map( A => n3459, Z => n1387);
   U438 : BUF_X1 port map( A => n3478, Z => n1354);
   U439 : BUF_X1 port map( A => n3481, Z => n1345);
   U440 : BUF_X1 port map( A => n3490, Z => n1321);
   U441 : BUF_X1 port map( A => n3509, Z => n1192);
   U442 : BUF_X1 port map( A => n3512, Z => n1183);
   U443 : BUF_X1 port map( A => n3515, Z => n1174);
   U444 : BUF_X1 port map( A => n4919, Z => n649);
   U445 : BUF_X1 port map( A => n3476, Z => n1361);
   U446 : BUF_X1 port map( A => n4950, Z => n487);
   U447 : BUF_X1 port map( A => n4981, Z => n69);
   U448 : BUF_X1 port map( A => n3538, Z => n781);
   U449 : BUF_X1 port map( A => n3507, Z => n1199);
   U450 : BUF_X1 port map( A => n4906, Z => n663);
   U451 : BUF_X1 port map( A => n4937, Z => n597);
   U452 : BUF_X1 port map( A => n4940, Z => n492);
   U453 : BUF_X1 port map( A => n4968, Z => n435);
   U454 : BUF_X1 port map( A => n4971, Z => n74);
   U455 : BUF_X1 port map( A => n4999, Z => n16);
   U456 : BUF_X1 port map( A => n5002, Z => n5);
   U457 : BUF_X1 port map( A => n3463, Z => n1375);
   U458 : BUF_X1 port map( A => n3494, Z => n1309);
   U459 : BUF_X1 port map( A => n3497, Z => n1300);
   U460 : BUF_X1 port map( A => n3525, Z => n1147);
   U461 : BUF_X1 port map( A => n3528, Z => n1138);
   U462 : BUF_X1 port map( A => n3556, Z => n729);
   U463 : BUF_X1 port map( A => n3559, Z => n720);
   U464 : BUF_X1 port map( A => n4906, Z => n662);
   U465 : BUF_X1 port map( A => n4937, Z => n596);
   U466 : BUF_X1 port map( A => n4940, Z => n491);
   U467 : BUF_X1 port map( A => n4968, Z => n434);
   U468 : BUF_X1 port map( A => n4971, Z => n73);
   U469 : BUF_X1 port map( A => n4999, Z => n15);
   U470 : BUF_X1 port map( A => n5002, Z => n4);
   U471 : BUF_X1 port map( A => n3463, Z => n1374);
   U472 : BUF_X1 port map( A => n3494, Z => n1308);
   U473 : BUF_X1 port map( A => n3497, Z => n1299);
   U474 : BUF_X1 port map( A => n3525, Z => n1146);
   U475 : BUF_X1 port map( A => n3528, Z => n1137);
   U476 : BUF_X1 port map( A => n3556, Z => n728);
   U477 : BUF_X1 port map( A => n3559, Z => n719);
   U478 : BUF_X1 port map( A => n4898, Z => n685);
   U479 : BUF_X1 port map( A => n4929, Z => n619);
   U480 : BUF_X1 port map( A => n4960, Z => n457);
   U481 : BUF_X1 port map( A => n4991, Z => n39);
   U482 : BUF_X1 port map( A => n3455, Z => n1397);
   U483 : BUF_X1 port map( A => n3486, Z => n1331);
   U484 : BUF_X1 port map( A => n3517, Z => n1169);
   U485 : BUF_X1 port map( A => n3548, Z => n751);
   U486 : BUF_X1 port map( A => n4904, Z => n670);
   U487 : BUF_X1 port map( A => n4907, Z => n661);
   U488 : BUF_X1 port map( A => n4935, Z => n604);
   U489 : BUF_X1 port map( A => n4938, Z => n595);
   U490 : BUF_X1 port map( A => n4966, Z => n442);
   U491 : BUF_X1 port map( A => n4969, Z => n433);
   U492 : BUF_X1 port map( A => n4997, Z => n24);
   U493 : BUF_X1 port map( A => n5000, Z => n14);
   U494 : BUF_X1 port map( A => n3461, Z => n1382);
   U495 : BUF_X1 port map( A => n3464, Z => n1373);
   U496 : BUF_X1 port map( A => n3492, Z => n1316);
   U497 : BUF_X1 port map( A => n3495, Z => n1307);
   U498 : BUF_X1 port map( A => n3523, Z => n1154);
   U499 : BUF_X1 port map( A => n3526, Z => n1145);
   U500 : BUF_X1 port map( A => n3554, Z => n736);
   U501 : BUF_X1 port map( A => n3557, Z => n727);
   U502 : BUF_X1 port map( A => n4899, Z => n682);
   U503 : BUF_X1 port map( A => n4930, Z => n616);
   U504 : BUF_X1 port map( A => n4961, Z => n454);
   U505 : BUF_X1 port map( A => n4992, Z => n36);
   U506 : BUF_X1 port map( A => n3456, Z => n1394);
   U507 : BUF_X1 port map( A => n3487, Z => n1328);
   U508 : BUF_X1 port map( A => n3518, Z => n1166);
   U509 : BUF_X1 port map( A => n3549, Z => n748);
   U510 : BUF_X1 port map( A => n3103, Z => n1744);
   U511 : BUF_X1 port map( A => n3103, Z => n1743);
   U512 : BUF_X1 port map( A => n3098, Z => n1747);
   U513 : BUF_X1 port map( A => n3098, Z => n1746);
   U514 : BUF_X1 port map( A => n3093, Z => n1750);
   U515 : BUF_X1 port map( A => n3093, Z => n1749);
   U516 : BUF_X1 port map( A => n3088, Z => n1753);
   U517 : BUF_X1 port map( A => n3088, Z => n1752);
   U518 : BUF_X1 port map( A => n3083, Z => n1756);
   U519 : BUF_X1 port map( A => n3083, Z => n1755);
   U520 : BUF_X1 port map( A => n3078, Z => n1759);
   U521 : BUF_X1 port map( A => n3078, Z => n1758);
   U522 : BUF_X1 port map( A => n3073, Z => n1762);
   U523 : BUF_X1 port map( A => n3073, Z => n1761);
   U524 : BUF_X1 port map( A => n3068, Z => n1765);
   U525 : BUF_X1 port map( A => n3068, Z => n1764);
   U526 : BUF_X1 port map( A => n3063, Z => n1768);
   U527 : BUF_X1 port map( A => n3063, Z => n1767);
   U528 : BUF_X1 port map( A => n3058, Z => n1771);
   U529 : BUF_X1 port map( A => n3058, Z => n1770);
   U530 : BUF_X1 port map( A => n3053, Z => n1774);
   U531 : BUF_X1 port map( A => n3053, Z => n1773);
   U532 : BUF_X1 port map( A => n3048, Z => n1777);
   U533 : BUF_X1 port map( A => n3048, Z => n1776);
   U534 : BUF_X1 port map( A => n3043, Z => n1780);
   U535 : BUF_X1 port map( A => n3043, Z => n1779);
   U536 : BUF_X1 port map( A => n3038, Z => n1783);
   U537 : BUF_X1 port map( A => n3038, Z => n1782);
   U538 : BUF_X1 port map( A => n3033, Z => n1786);
   U539 : BUF_X1 port map( A => n3033, Z => n1785);
   U540 : BUF_X1 port map( A => n2996, Z => n1789);
   U541 : BUF_X1 port map( A => n2996, Z => n1788);
   U542 : BUF_X1 port map( A => n3303, Z => n1504);
   U543 : BUF_X1 port map( A => n3303, Z => n1503);
   U544 : BUF_X1 port map( A => n3299, Z => n1507);
   U545 : BUF_X1 port map( A => n3299, Z => n1506);
   U546 : BUF_X1 port map( A => n3295, Z => n1510);
   U547 : BUF_X1 port map( A => n3295, Z => n1509);
   U548 : BUF_X1 port map( A => n3291, Z => n1513);
   U549 : BUF_X1 port map( A => n3291, Z => n1512);
   U550 : BUF_X1 port map( A => n3287, Z => n1516);
   U551 : BUF_X1 port map( A => n3287, Z => n1515);
   U552 : BUF_X1 port map( A => n3283, Z => n1519);
   U553 : BUF_X1 port map( A => n3283, Z => n1518);
   U554 : BUF_X1 port map( A => n3279, Z => n1522);
   U555 : BUF_X1 port map( A => n3279, Z => n1521);
   U556 : BUF_X1 port map( A => n3275, Z => n1525);
   U557 : BUF_X1 port map( A => n3275, Z => n1524);
   U558 : BUF_X1 port map( A => n3271, Z => n1528);
   U559 : BUF_X1 port map( A => n3271, Z => n1527);
   U560 : BUF_X1 port map( A => n3267, Z => n1531);
   U561 : BUF_X1 port map( A => n3267, Z => n1530);
   U562 : BUF_X1 port map( A => n3263, Z => n1534);
   U563 : BUF_X1 port map( A => n3263, Z => n1533);
   U564 : BUF_X1 port map( A => n3259, Z => n1537);
   U565 : BUF_X1 port map( A => n3259, Z => n1536);
   U566 : BUF_X1 port map( A => n3255, Z => n1540);
   U567 : BUF_X1 port map( A => n3255, Z => n1539);
   U568 : BUF_X1 port map( A => n3251, Z => n1543);
   U569 : BUF_X1 port map( A => n3251, Z => n1542);
   U570 : BUF_X1 port map( A => n3247, Z => n1546);
   U571 : BUF_X1 port map( A => n3247, Z => n1545);
   U572 : BUF_X1 port map( A => n3242, Z => n1549);
   U573 : BUF_X1 port map( A => n3242, Z => n1548);
   U574 : BUF_X1 port map( A => n3238, Z => n1648);
   U575 : BUF_X1 port map( A => n3238, Z => n1551);
   U576 : BUF_X1 port map( A => n3234, Z => n1651);
   U577 : BUF_X1 port map( A => n3234, Z => n1650);
   U578 : BUF_X1 port map( A => n3230, Z => n1654);
   U579 : BUF_X1 port map( A => n3230, Z => n1653);
   U580 : BUF_X1 port map( A => n3226, Z => n1657);
   U581 : BUF_X1 port map( A => n3226, Z => n1656);
   U582 : BUF_X1 port map( A => n3222, Z => n1660);
   U583 : BUF_X1 port map( A => n3222, Z => n1659);
   U584 : BUF_X1 port map( A => n3218, Z => n1663);
   U585 : BUF_X1 port map( A => n3218, Z => n1662);
   U586 : BUF_X1 port map( A => n3214, Z => n1666);
   U587 : BUF_X1 port map( A => n3214, Z => n1665);
   U588 : BUF_X1 port map( A => n3210, Z => n1669);
   U589 : BUF_X1 port map( A => n3210, Z => n1668);
   U590 : BUF_X1 port map( A => n3206, Z => n1672);
   U591 : BUF_X1 port map( A => n3206, Z => n1671);
   U592 : BUF_X1 port map( A => n3202, Z => n1675);
   U593 : BUF_X1 port map( A => n3202, Z => n1674);
   U594 : BUF_X1 port map( A => n3198, Z => n1678);
   U595 : BUF_X1 port map( A => n3198, Z => n1677);
   U596 : BUF_X1 port map( A => n3194, Z => n1681);
   U597 : BUF_X1 port map( A => n3194, Z => n1680);
   U598 : BUF_X1 port map( A => n3190, Z => n1684);
   U599 : BUF_X1 port map( A => n3190, Z => n1683);
   U600 : BUF_X1 port map( A => n3186, Z => n1687);
   U601 : BUF_X1 port map( A => n3186, Z => n1686);
   U602 : BUF_X1 port map( A => n3182, Z => n1690);
   U603 : BUF_X1 port map( A => n3182, Z => n1689);
   U604 : BUF_X1 port map( A => n3177, Z => n1693);
   U605 : BUF_X1 port map( A => n3177, Z => n1692);
   U606 : BUF_X1 port map( A => n3173, Z => n1696);
   U607 : BUF_X1 port map( A => n3173, Z => n1695);
   U608 : BUF_X1 port map( A => n3169, Z => n1699);
   U609 : BUF_X1 port map( A => n3169, Z => n1698);
   U610 : BUF_X1 port map( A => n3165, Z => n1702);
   U611 : BUF_X1 port map( A => n3165, Z => n1701);
   U612 : BUF_X1 port map( A => n3161, Z => n1705);
   U613 : BUF_X1 port map( A => n3161, Z => n1704);
   U614 : BUF_X1 port map( A => n3157, Z => n1708);
   U615 : BUF_X1 port map( A => n3157, Z => n1707);
   U616 : BUF_X1 port map( A => n3153, Z => n1711);
   U617 : BUF_X1 port map( A => n3153, Z => n1710);
   U618 : BUF_X1 port map( A => n3149, Z => n1714);
   U619 : BUF_X1 port map( A => n3149, Z => n1713);
   U620 : BUF_X1 port map( A => n3145, Z => n1717);
   U621 : BUF_X1 port map( A => n3145, Z => n1716);
   U622 : BUF_X1 port map( A => n3141, Z => n1720);
   U623 : BUF_X1 port map( A => n3141, Z => n1719);
   U624 : BUF_X1 port map( A => n3137, Z => n1723);
   U625 : BUF_X1 port map( A => n3137, Z => n1722);
   U626 : BUF_X1 port map( A => n3133, Z => n1726);
   U627 : BUF_X1 port map( A => n3133, Z => n1725);
   U628 : BUF_X1 port map( A => n3129, Z => n1729);
   U629 : BUF_X1 port map( A => n3129, Z => n1728);
   U630 : BUF_X1 port map( A => n3125, Z => n1732);
   U631 : BUF_X1 port map( A => n3125, Z => n1731);
   U632 : BUF_X1 port map( A => n3121, Z => n1735);
   U633 : BUF_X1 port map( A => n3121, Z => n1734);
   U634 : BUF_X1 port map( A => n3117, Z => n1738);
   U635 : BUF_X1 port map( A => n3117, Z => n1737);
   U636 : BUF_X1 port map( A => n3112, Z => n1741);
   U637 : BUF_X1 port map( A => n3112, Z => n1740);
   U638 : BUF_X1 port map( A => n3375, Z => n1456);
   U639 : BUF_X1 port map( A => n3375, Z => n1455);
   U640 : BUF_X1 port map( A => n3371, Z => n1459);
   U641 : BUF_X1 port map( A => n3371, Z => n1458);
   U642 : BUF_X1 port map( A => n3367, Z => n1462);
   U643 : BUF_X1 port map( A => n3367, Z => n1461);
   U644 : BUF_X1 port map( A => n3362, Z => n1465);
   U645 : BUF_X1 port map( A => n3362, Z => n1464);
   U646 : BUF_X1 port map( A => n3356, Z => n1468);
   U647 : BUF_X1 port map( A => n3356, Z => n1467);
   U648 : BUF_X1 port map( A => n3351, Z => n1471);
   U649 : BUF_X1 port map( A => n3351, Z => n1470);
   U650 : BUF_X1 port map( A => n3346, Z => n1474);
   U651 : BUF_X1 port map( A => n3346, Z => n1473);
   U652 : BUF_X1 port map( A => n3340, Z => n1477);
   U653 : BUF_X1 port map( A => n3340, Z => n1476);
   U654 : BUF_X1 port map( A => n3336, Z => n1480);
   U655 : BUF_X1 port map( A => n3336, Z => n1479);
   U656 : BUF_X1 port map( A => n3332, Z => n1483);
   U657 : BUF_X1 port map( A => n3332, Z => n1482);
   U658 : BUF_X1 port map( A => n3328, Z => n1486);
   U659 : BUF_X1 port map( A => n3328, Z => n1485);
   U660 : BUF_X1 port map( A => n3324, Z => n1489);
   U661 : BUF_X1 port map( A => n3324, Z => n1488);
   U662 : BUF_X1 port map( A => n3320, Z => n1492);
   U663 : BUF_X1 port map( A => n3320, Z => n1491);
   U664 : BUF_X1 port map( A => n3316, Z => n1495);
   U665 : BUF_X1 port map( A => n3316, Z => n1494);
   U666 : BUF_X1 port map( A => n3312, Z => n1498);
   U667 : BUF_X1 port map( A => n3312, Z => n1497);
   U668 : BUF_X1 port map( A => n3307, Z => n1501);
   U669 : BUF_X1 port map( A => n3307, Z => n1500);
   U670 : BUF_X1 port map( A => n3413, Z => n1432);
   U671 : BUF_X1 port map( A => n3413, Z => n1431);
   U672 : BUF_X1 port map( A => n3409, Z => n1435);
   U673 : BUF_X1 port map( A => n3409, Z => n1434);
   U674 : BUF_X1 port map( A => n3403, Z => n1438);
   U675 : BUF_X1 port map( A => n3403, Z => n1437);
   U676 : BUF_X1 port map( A => n3398, Z => n1441);
   U677 : BUF_X1 port map( A => n3398, Z => n1440);
   U678 : BUF_X1 port map( A => n3394, Z => n1444);
   U679 : BUF_X1 port map( A => n3394, Z => n1443);
   U680 : BUF_X1 port map( A => n3390, Z => n1447);
   U681 : BUF_X1 port map( A => n3390, Z => n1446);
   U682 : BUF_X1 port map( A => n3386, Z => n1450);
   U683 : BUF_X1 port map( A => n3386, Z => n1449);
   U684 : BUF_X1 port map( A => n3380, Z => n1453);
   U685 : BUF_X1 port map( A => n3380, Z => n1452);
   U686 : BUF_X1 port map( A => n4891, Z => n706);
   U687 : BUF_X1 port map( A => n3448, Z => n1418);
   U688 : BUF_X1 port map( A => n4990, Z => n42);
   U689 : BUF_X1 port map( A => n4996, Z => n27);
   U690 : BUF_X1 port map( A => n3547, Z => n754);
   U691 : BUF_X1 port map( A => n3553, Z => n739);
   U692 : BUF_X1 port map( A => n4894, Z => n697);
   U693 : BUF_X1 port map( A => n4984, Z => n60);
   U694 : BUF_X1 port map( A => n3451, Z => n1409);
   U695 : BUF_X1 port map( A => n3541, Z => n772);
   U696 : BUF_X1 port map( A => n4897, Z => n688);
   U697 : BUF_X1 port map( A => n4903, Z => n673);
   U698 : BUF_X1 port map( A => n4922, Z => n640);
   U699 : BUF_X1 port map( A => n4925, Z => n631);
   U700 : BUF_X1 port map( A => n4928, Z => n622);
   U701 : BUF_X1 port map( A => n4934, Z => n607);
   U702 : BUF_X1 port map( A => n4953, Z => n478);
   U703 : BUF_X1 port map( A => n4956, Z => n469);
   U704 : BUF_X1 port map( A => n4959, Z => n460);
   U705 : BUF_X1 port map( A => n4965, Z => n445);
   U706 : BUF_X1 port map( A => n4987, Z => n51);
   U707 : BUF_X1 port map( A => n3454, Z => n1400);
   U708 : BUF_X1 port map( A => n3460, Z => n1385);
   U709 : BUF_X1 port map( A => n3479, Z => n1352);
   U710 : BUF_X1 port map( A => n3482, Z => n1343);
   U711 : BUF_X1 port map( A => n3485, Z => n1334);
   U712 : BUF_X1 port map( A => n3491, Z => n1319);
   U713 : BUF_X1 port map( A => n3510, Z => n1190);
   U714 : BUF_X1 port map( A => n3513, Z => n1181);
   U715 : BUF_X1 port map( A => n3516, Z => n1172);
   U716 : BUF_X1 port map( A => n3522, Z => n1157);
   U717 : BUF_X1 port map( A => n3544, Z => n763);
   U718 : BUF_X1 port map( A => n4905, Z => n667);
   U719 : BUF_X1 port map( A => n4908, Z => n658);
   U720 : BUF_X1 port map( A => n4936, Z => n601);
   U721 : BUF_X1 port map( A => n4939, Z => n592);
   U722 : BUF_X1 port map( A => n4967, Z => n439);
   U723 : BUF_X1 port map( A => n4970, Z => n78);
   U724 : BUF_X1 port map( A => n4998, Z => n21);
   U725 : BUF_X1 port map( A => n5001, Z => n10);
   U726 : BUF_X1 port map( A => n3462, Z => n1379);
   U727 : BUF_X1 port map( A => n3465, Z => n1370);
   U728 : BUF_X1 port map( A => n3493, Z => n1313);
   U729 : BUF_X1 port map( A => n3496, Z => n1304);
   U730 : BUF_X1 port map( A => n3524, Z => n1151);
   U731 : BUF_X1 port map( A => n3527, Z => n1142);
   U732 : BUF_X1 port map( A => n3555, Z => n733);
   U733 : BUF_X1 port map( A => n3558, Z => n724);
   U734 : BUF_X1 port map( A => n4889, Z => n712);
   U735 : BUF_X1 port map( A => n3446, Z => n1424);
   U736 : BUF_X1 port map( A => n4985, Z => n57);
   U737 : BUF_X1 port map( A => n4988, Z => n48);
   U738 : BUF_X1 port map( A => n3542, Z => n769);
   U739 : BUF_X1 port map( A => n3545, Z => n760);
   U740 : BUF_X1 port map( A => n4892, Z => n703);
   U741 : BUF_X1 port map( A => n3449, Z => n1415);
   U742 : BUF_X1 port map( A => n4932, Z => n613);
   U743 : BUF_X1 port map( A => n3489, Z => n1325);
   U744 : BUF_X1 port map( A => n4895, Z => n694);
   U745 : BUF_X1 port map( A => n4901, Z => n679);
   U746 : BUF_X1 port map( A => n4920, Z => n646);
   U747 : BUF_X1 port map( A => n4923, Z => n637);
   U748 : BUF_X1 port map( A => n4926, Z => n628);
   U749 : BUF_X1 port map( A => n4951, Z => n484);
   U750 : BUF_X1 port map( A => n4954, Z => n475);
   U751 : BUF_X1 port map( A => n4963, Z => n451);
   U752 : BUF_X1 port map( A => n4982, Z => n66);
   U753 : BUF_X1 port map( A => n3539, Z => n778);
   U754 : BUF_X1 port map( A => n4994, Z => n33);
   U755 : BUF_X1 port map( A => n3452, Z => n1406);
   U756 : BUF_X1 port map( A => n3458, Z => n1391);
   U757 : BUF_X1 port map( A => n3477, Z => n1358);
   U758 : BUF_X1 port map( A => n3480, Z => n1349);
   U759 : BUF_X1 port map( A => n3483, Z => n1340);
   U760 : BUF_X1 port map( A => n3508, Z => n1196);
   U761 : BUF_X1 port map( A => n3511, Z => n1187);
   U762 : BUF_X1 port map( A => n3520, Z => n1163);
   U763 : BUF_X1 port map( A => n3551, Z => n745);
   U764 : BUF_X1 port map( A => n4986, Z => n54);
   U765 : BUF_X1 port map( A => n4989, Z => n45);
   U766 : BUF_X1 port map( A => n3543, Z => n766);
   U767 : BUF_X1 port map( A => n3546, Z => n757);
   U768 : BUF_X1 port map( A => n4893, Z => n700);
   U769 : BUF_X1 port map( A => n4983, Z => n63);
   U770 : BUF_X1 port map( A => n3450, Z => n1412);
   U771 : BUF_X1 port map( A => n3540, Z => n775);
   U772 : BUF_X1 port map( A => n4890, Z => n709);
   U773 : BUF_X1 port map( A => n3447, Z => n1421);
   U774 : BUF_X1 port map( A => n4896, Z => n691);
   U775 : BUF_X1 port map( A => n4902, Z => n676);
   U776 : BUF_X1 port map( A => n4921, Z => n643);
   U777 : BUF_X1 port map( A => n4924, Z => n634);
   U778 : BUF_X1 port map( A => n4933, Z => n610);
   U779 : BUF_X1 port map( A => n4952, Z => n481);
   U780 : BUF_X1 port map( A => n4955, Z => n472);
   U781 : BUF_X1 port map( A => n4958, Z => n463);
   U782 : BUF_X1 port map( A => n3453, Z => n1403);
   U783 : BUF_X1 port map( A => n3459, Z => n1388);
   U784 : BUF_X1 port map( A => n3478, Z => n1355);
   U785 : BUF_X1 port map( A => n3481, Z => n1346);
   U786 : BUF_X1 port map( A => n3490, Z => n1322);
   U787 : BUF_X1 port map( A => n3509, Z => n1193);
   U788 : BUF_X1 port map( A => n3512, Z => n1184);
   U789 : BUF_X1 port map( A => n3515, Z => n1175);
   U790 : BUF_X1 port map( A => n5002, Z => n6);
   U791 : BUF_X1 port map( A => n3559, Z => n721);
   U792 : BUF_X1 port map( A => n4906, Z => n664);
   U793 : BUF_X1 port map( A => n4937, Z => n598);
   U794 : BUF_X1 port map( A => n4940, Z => n493);
   U795 : BUF_X1 port map( A => n4968, Z => n436);
   U796 : BUF_X1 port map( A => n4971, Z => n75);
   U797 : BUF_X1 port map( A => n4999, Z => n18);
   U798 : BUF_X1 port map( A => n3463, Z => n1376);
   U799 : BUF_X1 port map( A => n3494, Z => n1310);
   U800 : BUF_X1 port map( A => n3497, Z => n1301);
   U801 : BUF_X1 port map( A => n3525, Z => n1148);
   U802 : BUF_X1 port map( A => n3528, Z => n1139);
   U803 : BUF_X1 port map( A => n3556, Z => n730);
   U804 : NAND2_X1 port map( A1 => n6247, A2 => n6312, ZN => n4995);
   U805 : NAND2_X1 port map( A1 => n4804, A2 => n4869, ZN => n3552);
   U806 : BUF_X1 port map( A => n3103, Z => n1745);
   U807 : BUF_X1 port map( A => n3098, Z => n1748);
   U808 : BUF_X1 port map( A => n3093, Z => n1751);
   U809 : BUF_X1 port map( A => n3088, Z => n1754);
   U810 : BUF_X1 port map( A => n3083, Z => n1757);
   U811 : BUF_X1 port map( A => n3078, Z => n1760);
   U812 : BUF_X1 port map( A => n3073, Z => n1763);
   U813 : BUF_X1 port map( A => n3068, Z => n1766);
   U814 : BUF_X1 port map( A => n3063, Z => n1769);
   U815 : BUF_X1 port map( A => n3058, Z => n1772);
   U816 : BUF_X1 port map( A => n3053, Z => n1775);
   U817 : BUF_X1 port map( A => n3048, Z => n1778);
   U818 : BUF_X1 port map( A => n3043, Z => n1781);
   U819 : BUF_X1 port map( A => n3038, Z => n1784);
   U820 : BUF_X1 port map( A => n3033, Z => n1787);
   U821 : BUF_X1 port map( A => n2996, Z => n1790);
   U822 : BUF_X1 port map( A => n3303, Z => n1505);
   U823 : BUF_X1 port map( A => n3299, Z => n1508);
   U824 : BUF_X1 port map( A => n3295, Z => n1511);
   U825 : BUF_X1 port map( A => n3291, Z => n1514);
   U826 : BUF_X1 port map( A => n3287, Z => n1517);
   U827 : BUF_X1 port map( A => n3283, Z => n1520);
   U828 : BUF_X1 port map( A => n3279, Z => n1523);
   U829 : BUF_X1 port map( A => n3275, Z => n1526);
   U830 : BUF_X1 port map( A => n3271, Z => n1529);
   U831 : BUF_X1 port map( A => n3267, Z => n1532);
   U832 : BUF_X1 port map( A => n3263, Z => n1535);
   U833 : BUF_X1 port map( A => n3259, Z => n1538);
   U834 : BUF_X1 port map( A => n3255, Z => n1541);
   U835 : BUF_X1 port map( A => n3251, Z => n1544);
   U836 : BUF_X1 port map( A => n3247, Z => n1547);
   U837 : BUF_X1 port map( A => n3242, Z => n1550);
   U838 : BUF_X1 port map( A => n3238, Z => n1649);
   U839 : BUF_X1 port map( A => n3234, Z => n1652);
   U840 : BUF_X1 port map( A => n3230, Z => n1655);
   U841 : BUF_X1 port map( A => n3226, Z => n1658);
   U842 : BUF_X1 port map( A => n3222, Z => n1661);
   U843 : BUF_X1 port map( A => n3218, Z => n1664);
   U844 : BUF_X1 port map( A => n3214, Z => n1667);
   U845 : BUF_X1 port map( A => n3210, Z => n1670);
   U846 : BUF_X1 port map( A => n3206, Z => n1673);
   U847 : BUF_X1 port map( A => n3202, Z => n1676);
   U848 : BUF_X1 port map( A => n3198, Z => n1679);
   U849 : BUF_X1 port map( A => n3194, Z => n1682);
   U850 : BUF_X1 port map( A => n3190, Z => n1685);
   U851 : BUF_X1 port map( A => n3186, Z => n1688);
   U852 : BUF_X1 port map( A => n3182, Z => n1691);
   U853 : BUF_X1 port map( A => n3177, Z => n1694);
   U854 : BUF_X1 port map( A => n3173, Z => n1697);
   U855 : BUF_X1 port map( A => n3169, Z => n1700);
   U856 : BUF_X1 port map( A => n3165, Z => n1703);
   U857 : BUF_X1 port map( A => n3161, Z => n1706);
   U858 : BUF_X1 port map( A => n3157, Z => n1709);
   U859 : BUF_X1 port map( A => n3153, Z => n1712);
   U860 : BUF_X1 port map( A => n3149, Z => n1715);
   U861 : BUF_X1 port map( A => n3145, Z => n1718);
   U862 : BUF_X1 port map( A => n3141, Z => n1721);
   U863 : BUF_X1 port map( A => n3137, Z => n1724);
   U864 : BUF_X1 port map( A => n3133, Z => n1727);
   U865 : BUF_X1 port map( A => n3129, Z => n1730);
   U866 : BUF_X1 port map( A => n3125, Z => n1733);
   U867 : BUF_X1 port map( A => n3121, Z => n1736);
   U868 : BUF_X1 port map( A => n3117, Z => n1739);
   U869 : BUF_X1 port map( A => n3112, Z => n1742);
   U870 : BUF_X1 port map( A => n3375, Z => n1457);
   U871 : BUF_X1 port map( A => n3371, Z => n1460);
   U872 : BUF_X1 port map( A => n3367, Z => n1463);
   U873 : BUF_X1 port map( A => n3362, Z => n1466);
   U874 : BUF_X1 port map( A => n3356, Z => n1469);
   U875 : BUF_X1 port map( A => n3351, Z => n1472);
   U876 : BUF_X1 port map( A => n3346, Z => n1475);
   U877 : BUF_X1 port map( A => n3340, Z => n1478);
   U878 : BUF_X1 port map( A => n3336, Z => n1481);
   U879 : BUF_X1 port map( A => n3332, Z => n1484);
   U880 : BUF_X1 port map( A => n3328, Z => n1487);
   U881 : BUF_X1 port map( A => n3324, Z => n1490);
   U882 : BUF_X1 port map( A => n3320, Z => n1493);
   U883 : BUF_X1 port map( A => n3316, Z => n1496);
   U884 : BUF_X1 port map( A => n3312, Z => n1499);
   U885 : BUF_X1 port map( A => n3307, Z => n1502);
   U886 : BUF_X1 port map( A => n3413, Z => n1433);
   U887 : BUF_X1 port map( A => n3409, Z => n1436);
   U888 : BUF_X1 port map( A => n3403, Z => n1439);
   U889 : BUF_X1 port map( A => n3398, Z => n1442);
   U890 : BUF_X1 port map( A => n3394, Z => n1445);
   U891 : BUF_X1 port map( A => n3390, Z => n1448);
   U892 : BUF_X1 port map( A => n3386, Z => n1451);
   U893 : BUF_X1 port map( A => n3380, Z => n1454);
   U894 : NAND2_X1 port map( A1 => n6248, A2 => n6247, ZN => n4887);
   U895 : NAND2_X1 port map( A1 => n6246, A2 => n6247, ZN => n4888);
   U896 : NAND2_X1 port map( A1 => n6281, A2 => n6247, ZN => n4927);
   U897 : NAND2_X1 port map( A1 => n6298, A2 => n6247, ZN => n4957);
   U898 : NAND2_X1 port map( A1 => n6300, A2 => n6247, ZN => n4964);
   U899 : NAND2_X1 port map( A1 => n4805, A2 => n4804, ZN => n3444);
   U900 : NAND2_X1 port map( A1 => n4803, A2 => n4804, ZN => n3445);
   U901 : NAND2_X1 port map( A1 => n4838, A2 => n4804, ZN => n3484);
   U902 : NAND2_X1 port map( A1 => n4855, A2 => n4804, ZN => n3514);
   U903 : NAND2_X1 port map( A1 => n4857, A2 => n4804, ZN => n3521);
   U904 : AND2_X1 port map( A1 => n6268, A2 => n6247, ZN => n4909);
   U905 : AND2_X1 port map( A1 => n4825, A2 => n4804, ZN => n3466);
   U906 : INV_X1 port map( A => n2955, ZN => n3363);
   U907 : NOR2_X1 port map( A1 => n3372, A2 => n3373, ZN => n3343);
   U908 : NOR2_X1 port map( A1 => n3369, A2 => n3370, ZN => n3383);
   U909 : NAND2_X1 port map( A1 => n3400, A2 => n3358, ZN => n3065);
   U910 : NAND2_X1 port map( A1 => n3400, A2 => n3353, ZN => n3060);
   U911 : NAND2_X1 port map( A1 => n3400, A2 => n3348, ZN => n3055);
   U912 : NAND2_X1 port map( A1 => n3400, A2 => n3343, ZN => n3050);
   U913 : NAND2_X1 port map( A1 => n3358, A2 => n3383, ZN => n3045);
   U914 : NAND2_X1 port map( A1 => n3353, A2 => n3383, ZN => n3040);
   U915 : NAND2_X1 port map( A1 => n3348, A2 => n3383, ZN => n3035);
   U916 : NOR2_X1 port map( A1 => n3029, A2 => n3105, ZN => n3103);
   U917 : NOR2_X1 port map( A1 => n3029, A2 => n3100, ZN => n3098);
   U918 : NOR2_X1 port map( A1 => n3029, A2 => n3095, ZN => n3093);
   U919 : NOR2_X1 port map( A1 => n3029, A2 => n3090, ZN => n3088);
   U920 : NOR2_X1 port map( A1 => n3029, A2 => n3085, ZN => n3083);
   U921 : NOR2_X1 port map( A1 => n3029, A2 => n3080, ZN => n3078);
   U922 : NOR2_X1 port map( A1 => n3029, A2 => n3075, ZN => n3073);
   U923 : NOR2_X1 port map( A1 => n3029, A2 => n3070, ZN => n3068);
   U924 : NOR2_X1 port map( A1 => n3029, A2 => n3065, ZN => n3063);
   U925 : NOR2_X1 port map( A1 => n3029, A2 => n3060, ZN => n3058);
   U926 : NOR2_X1 port map( A1 => n3029, A2 => n3055, ZN => n3053);
   U927 : NOR2_X1 port map( A1 => n3029, A2 => n3050, ZN => n3048);
   U928 : NOR2_X1 port map( A1 => n3029, A2 => n3045, ZN => n3043);
   U929 : NOR2_X1 port map( A1 => n3029, A2 => n3040, ZN => n3038);
   U930 : NOR2_X1 port map( A1 => n3029, A2 => n3035, ZN => n3033);
   U931 : NOR2_X1 port map( A1 => n3029, A2 => n3030, ZN => n2996);
   U932 : NAND2_X1 port map( A1 => n3364, A2 => n3358, ZN => n3105);
   U933 : NAND2_X1 port map( A1 => n3364, A2 => n3353, ZN => n3100);
   U934 : NAND2_X1 port map( A1 => n3342, A2 => n3358, ZN => n3085);
   U935 : NAND2_X1 port map( A1 => n3342, A2 => n3353, ZN => n3080);
   U936 : NAND2_X1 port map( A1 => n3364, A2 => n3348, ZN => n3095);
   U937 : NAND2_X1 port map( A1 => n3342, A2 => n3348, ZN => n3075);
   U938 : NAND2_X1 port map( A1 => n3364, A2 => n3343, ZN => n3090);
   U939 : NAND2_X1 port map( A1 => n3342, A2 => n3343, ZN => n3070);
   U940 : NOR2_X1 port map( A1 => n3105, A2 => n3244, ZN => n3303);
   U941 : NOR2_X1 port map( A1 => n3100, A2 => n3244, ZN => n3299);
   U942 : NOR2_X1 port map( A1 => n3095, A2 => n3244, ZN => n3295);
   U943 : NOR2_X1 port map( A1 => n3090, A2 => n3244, ZN => n3291);
   U944 : NOR2_X1 port map( A1 => n3085, A2 => n3244, ZN => n3287);
   U945 : NOR2_X1 port map( A1 => n3080, A2 => n3244, ZN => n3283);
   U946 : NOR2_X1 port map( A1 => n3075, A2 => n3244, ZN => n3279);
   U947 : NOR2_X1 port map( A1 => n3070, A2 => n3244, ZN => n3275);
   U948 : NOR2_X1 port map( A1 => n3065, A2 => n3244, ZN => n3271);
   U949 : NOR2_X1 port map( A1 => n3060, A2 => n3244, ZN => n3267);
   U950 : NOR2_X1 port map( A1 => n3055, A2 => n3244, ZN => n3263);
   U951 : NOR2_X1 port map( A1 => n3050, A2 => n3244, ZN => n3259);
   U952 : NOR2_X1 port map( A1 => n3045, A2 => n3244, ZN => n3255);
   U953 : NOR2_X1 port map( A1 => n3040, A2 => n3244, ZN => n3251);
   U954 : NOR2_X1 port map( A1 => n3035, A2 => n3244, ZN => n3247);
   U955 : NOR2_X1 port map( A1 => n3030, A2 => n3244, ZN => n3242);
   U956 : NOR2_X1 port map( A1 => n3105, A2 => n3179, ZN => n3238);
   U957 : NOR2_X1 port map( A1 => n3100, A2 => n3179, ZN => n3234);
   U958 : NOR2_X1 port map( A1 => n3095, A2 => n3179, ZN => n3230);
   U959 : NOR2_X1 port map( A1 => n3090, A2 => n3179, ZN => n3226);
   U960 : NOR2_X1 port map( A1 => n3085, A2 => n3179, ZN => n3222);
   U961 : NOR2_X1 port map( A1 => n3080, A2 => n3179, ZN => n3218);
   U962 : NOR2_X1 port map( A1 => n3075, A2 => n3179, ZN => n3214);
   U963 : NOR2_X1 port map( A1 => n3070, A2 => n3179, ZN => n3210);
   U964 : NOR2_X1 port map( A1 => n3065, A2 => n3179, ZN => n3206);
   U965 : NOR2_X1 port map( A1 => n3060, A2 => n3179, ZN => n3202);
   U966 : NOR2_X1 port map( A1 => n3055, A2 => n3179, ZN => n3198);
   U967 : NOR2_X1 port map( A1 => n3050, A2 => n3179, ZN => n3194);
   U968 : NOR2_X1 port map( A1 => n3045, A2 => n3179, ZN => n3190);
   U969 : NOR2_X1 port map( A1 => n3040, A2 => n3179, ZN => n3186);
   U970 : NOR2_X1 port map( A1 => n3035, A2 => n3179, ZN => n3182);
   U971 : NOR2_X1 port map( A1 => n3030, A2 => n3179, ZN => n3177);
   U972 : NOR2_X1 port map( A1 => n3105, A2 => n3114, ZN => n3173);
   U973 : NOR2_X1 port map( A1 => n3100, A2 => n3114, ZN => n3169);
   U974 : NOR2_X1 port map( A1 => n3095, A2 => n3114, ZN => n3165);
   U975 : NOR2_X1 port map( A1 => n3090, A2 => n3114, ZN => n3161);
   U976 : NOR2_X1 port map( A1 => n3085, A2 => n3114, ZN => n3157);
   U977 : NOR2_X1 port map( A1 => n3080, A2 => n3114, ZN => n3153);
   U978 : NOR2_X1 port map( A1 => n3075, A2 => n3114, ZN => n3149);
   U979 : NOR2_X1 port map( A1 => n3070, A2 => n3114, ZN => n3145);
   U980 : NOR2_X1 port map( A1 => n3065, A2 => n3114, ZN => n3141);
   U981 : NOR2_X1 port map( A1 => n3060, A2 => n3114, ZN => n3137);
   U982 : NOR2_X1 port map( A1 => n3055, A2 => n3114, ZN => n3133);
   U983 : NOR2_X1 port map( A1 => n3050, A2 => n3114, ZN => n3129);
   U984 : NOR2_X1 port map( A1 => n3045, A2 => n3114, ZN => n3125);
   U985 : NOR2_X1 port map( A1 => n3040, A2 => n3114, ZN => n3121);
   U986 : NOR2_X1 port map( A1 => n3035, A2 => n3114, ZN => n3117);
   U987 : NOR2_X1 port map( A1 => n3030, A2 => n3114, ZN => n3112);
   U988 : NOR2_X1 port map( A1 => n3105, A2 => n3309, ZN => n3375);
   U989 : NOR2_X1 port map( A1 => n3100, A2 => n3309, ZN => n3371);
   U990 : NOR2_X1 port map( A1 => n3095, A2 => n3309, ZN => n3367);
   U991 : NOR2_X1 port map( A1 => n3090, A2 => n3309, ZN => n3362);
   U992 : NOR2_X1 port map( A1 => n3085, A2 => n3309, ZN => n3356);
   U993 : NOR2_X1 port map( A1 => n3080, A2 => n3309, ZN => n3351);
   U994 : NOR2_X1 port map( A1 => n3075, A2 => n3309, ZN => n3346);
   U995 : NOR2_X1 port map( A1 => n3070, A2 => n3309, ZN => n3340);
   U996 : NOR2_X1 port map( A1 => n3065, A2 => n3309, ZN => n3336);
   U997 : NOR2_X1 port map( A1 => n3060, A2 => n3309, ZN => n3332);
   U998 : NOR2_X1 port map( A1 => n3055, A2 => n3309, ZN => n3328);
   U999 : NOR2_X1 port map( A1 => n3050, A2 => n3309, ZN => n3324);
   U1000 : NOR2_X1 port map( A1 => n3045, A2 => n3309, ZN => n3320);
   U1001 : NOR2_X1 port map( A1 => n3040, A2 => n3309, ZN => n3316);
   U1002 : NOR2_X1 port map( A1 => n3035, A2 => n3309, ZN => n3312);
   U1003 : NOR2_X1 port map( A1 => n3030, A2 => n3309, ZN => n3307);
   U1004 : AND2_X1 port map( A1 => n6309, A2 => n6251, ZN => n6260);
   U1005 : AND2_X1 port map( A1 => n4866, A2 => n4808, ZN => n4817);
   U1006 : NOR2_X1 port map( A1 => n3065, A2 => n3382, ZN => n3413);
   U1007 : NOR2_X1 port map( A1 => n3060, A2 => n3382, ZN => n3409);
   U1008 : NOR2_X1 port map( A1 => n3055, A2 => n3382, ZN => n3403);
   U1009 : NOR2_X1 port map( A1 => n3050, A2 => n3382, ZN => n3398);
   U1010 : NOR2_X1 port map( A1 => n3045, A2 => n3382, ZN => n3394);
   U1011 : NOR2_X1 port map( A1 => n3040, A2 => n3382, ZN => n3390);
   U1012 : NOR2_X1 port map( A1 => n3035, A2 => n3382, ZN => n3386);
   U1013 : NOR2_X1 port map( A1 => n3030, A2 => n3382, ZN => n3380);
   U1014 : AND2_X1 port map( A1 => n6310, A2 => n6251, ZN => n6261);
   U1015 : AND2_X1 port map( A1 => n4867, A2 => n4808, ZN => n4818);
   U1016 : AND2_X1 port map( A1 => n6310, A2 => n6249, ZN => n6256);
   U1017 : AND2_X1 port map( A1 => n4867, A2 => n4806, ZN => n4813);
   U1018 : AND2_X1 port map( A1 => n6310, A2 => n6247, ZN => n6255);
   U1019 : AND2_X1 port map( A1 => n6309, A2 => n6247, ZN => n6257);
   U1020 : AND2_X1 port map( A1 => n4867, A2 => n4804, ZN => n4812);
   U1021 : AND2_X1 port map( A1 => n4866, A2 => n4804, ZN => n4814);
   U1022 : AND2_X1 port map( A1 => n6309, A2 => n6250, ZN => n6259);
   U1023 : AND2_X1 port map( A1 => n4866, A2 => n4807, ZN => n4816);
   U1024 : AND2_X1 port map( A1 => n6309, A2 => n6249, ZN => n6262);
   U1025 : AND2_X1 port map( A1 => n4866, A2 => n4806, ZN => n4819);
   U1026 : AND2_X1 port map( A1 => n6310, A2 => n6250, ZN => n6263);
   U1027 : AND2_X1 port map( A1 => n4867, A2 => n4807, ZN => n4820);
   U1028 : NAND2_X1 port map( A1 => n6296, A2 => n6257, ZN => n4953);
   U1029 : NAND2_X1 port map( A1 => n6296, A2 => n6256, ZN => n4951);
   U1030 : NAND2_X1 port map( A1 => n6296, A2 => n6262, ZN => n4952);
   U1031 : NAND2_X1 port map( A1 => n6296, A2 => n6263, ZN => n4956);
   U1032 : NAND2_X1 port map( A1 => n6296, A2 => n6259, ZN => n4954);
   U1033 : NAND2_X1 port map( A1 => n6296, A2 => n6261, ZN => n4955);
   U1034 : NAND2_X1 port map( A1 => n6296, A2 => n6260, ZN => n4959);
   U1035 : NAND2_X1 port map( A1 => n6296, A2 => n6287, ZN => n4949);
   U1036 : NAND2_X1 port map( A1 => n6296, A2 => n6255, ZN => n4950);
   U1037 : NAND2_X1 port map( A1 => n4853, A2 => n4814, ZN => n3510);
   U1038 : NAND2_X1 port map( A1 => n4853, A2 => n4813, ZN => n3508);
   U1039 : NAND2_X1 port map( A1 => n4853, A2 => n4819, ZN => n3509);
   U1040 : NAND2_X1 port map( A1 => n4853, A2 => n4820, ZN => n3513);
   U1041 : NAND2_X1 port map( A1 => n4853, A2 => n4816, ZN => n3511);
   U1042 : NAND2_X1 port map( A1 => n4853, A2 => n4818, ZN => n3512);
   U1043 : NAND2_X1 port map( A1 => n4853, A2 => n4817, ZN => n3516);
   U1044 : NAND2_X1 port map( A1 => n4853, A2 => n4844, ZN => n3506);
   U1045 : NAND2_X1 port map( A1 => n4853, A2 => n4812, ZN => n3507);
   U1046 : NAND2_X1 port map( A1 => n6248, A2 => n6249, ZN => n4891);
   U1047 : NAND2_X1 port map( A1 => n6246, A2 => n6249, ZN => n4889);
   U1048 : NAND2_X1 port map( A1 => n6298, A2 => n6249, ZN => n4980);
   U1049 : NAND2_X1 port map( A1 => n4805, A2 => n4806, ZN => n3448);
   U1050 : NAND2_X1 port map( A1 => n4803, A2 => n4806, ZN => n3446);
   U1051 : NAND2_X1 port map( A1 => n4855, A2 => n4806, ZN => n3537);
   U1052 : BUF_X1 port map( A => n1797, Z => n1800);
   U1053 : BUF_X1 port map( A => n1808, Z => n1811);
   U1054 : BUF_X1 port map( A => n1819, Z => n1822);
   U1055 : BUF_X1 port map( A => n1830, Z => n1833);
   U1056 : BUF_X1 port map( A => n2545, Z => n2548);
   U1057 : BUF_X1 port map( A => n2556, Z => n2559);
   U1058 : BUF_X1 port map( A => n2567, Z => n2570);
   U1059 : BUF_X1 port map( A => n2578, Z => n2581);
   U1060 : BUF_X1 port map( A => n2589, Z => n2592);
   U1061 : BUF_X1 port map( A => n2600, Z => n2603);
   U1062 : BUF_X1 port map( A => n2707, Z => n2710);
   U1063 : BUF_X1 port map( A => n2718, Z => n2721);
   U1064 : BUF_X1 port map( A => n2729, Z => n2732);
   U1065 : BUF_X1 port map( A => n2740, Z => n2743);
   U1066 : BUF_X1 port map( A => n2751, Z => n2754);
   U1067 : BUF_X1 port map( A => n2762, Z => n2765);
   U1068 : BUF_X1 port map( A => n2773, Z => n2776);
   U1069 : BUF_X1 port map( A => n2784, Z => n2787);
   U1070 : BUF_X1 port map( A => n2795, Z => n2798);
   U1071 : BUF_X1 port map( A => n2806, Z => n2809);
   U1072 : BUF_X1 port map( A => n2817, Z => n2820);
   U1073 : BUF_X1 port map( A => n2828, Z => n2831);
   U1074 : BUF_X1 port map( A => n2839, Z => n2842);
   U1075 : BUF_X1 port map( A => n2850, Z => n2853);
   U1076 : BUF_X1 port map( A => n2861, Z => n2864);
   U1077 : BUF_X1 port map( A => n2872, Z => n2875);
   U1078 : BUF_X1 port map( A => n2883, Z => n2886);
   U1079 : BUF_X1 port map( A => n2894, Z => n2897);
   U1080 : BUF_X1 port map( A => n2906, Z => n2909);
   U1081 : BUF_X1 port map( A => n2922, Z => n2925);
   U1082 : BUF_X1 port map( A => n2933, Z => n2936);
   U1083 : BUF_X1 port map( A => n2944, Z => n2947);
   U1084 : BUF_X1 port map( A => n1797, Z => n1801);
   U1085 : BUF_X1 port map( A => n1808, Z => n1812);
   U1086 : BUF_X1 port map( A => n1819, Z => n1823);
   U1087 : BUF_X1 port map( A => n1830, Z => n1834);
   U1088 : BUF_X1 port map( A => n2545, Z => n2549);
   U1089 : BUF_X1 port map( A => n2556, Z => n2560);
   U1090 : BUF_X1 port map( A => n2567, Z => n2571);
   U1091 : BUF_X1 port map( A => n2578, Z => n2582);
   U1092 : BUF_X1 port map( A => n2589, Z => n2593);
   U1093 : BUF_X1 port map( A => n2600, Z => n2604);
   U1094 : BUF_X1 port map( A => n2707, Z => n2711);
   U1095 : BUF_X1 port map( A => n2718, Z => n2722);
   U1096 : BUF_X1 port map( A => n2729, Z => n2733);
   U1097 : BUF_X1 port map( A => n2740, Z => n2744);
   U1098 : BUF_X1 port map( A => n2751, Z => n2755);
   U1099 : BUF_X1 port map( A => n2762, Z => n2766);
   U1100 : BUF_X1 port map( A => n2773, Z => n2777);
   U1101 : BUF_X1 port map( A => n2784, Z => n2788);
   U1102 : BUF_X1 port map( A => n2795, Z => n2799);
   U1103 : BUF_X1 port map( A => n2806, Z => n2810);
   U1104 : BUF_X1 port map( A => n2817, Z => n2821);
   U1105 : BUF_X1 port map( A => n2828, Z => n2832);
   U1106 : BUF_X1 port map( A => n2839, Z => n2843);
   U1107 : BUF_X1 port map( A => n2850, Z => n2854);
   U1108 : BUF_X1 port map( A => n2861, Z => n2865);
   U1109 : BUF_X1 port map( A => n2872, Z => n2876);
   U1110 : BUF_X1 port map( A => n2883, Z => n2887);
   U1111 : BUF_X1 port map( A => n2894, Z => n2899);
   U1112 : BUF_X1 port map( A => n2906, Z => n2910);
   U1113 : BUF_X1 port map( A => n2922, Z => n2926);
   U1114 : BUF_X1 port map( A => n2933, Z => n2937);
   U1115 : BUF_X1 port map( A => n2944, Z => n2948);
   U1116 : BUF_X1 port map( A => n1797, Z => n1802);
   U1117 : BUF_X1 port map( A => n1808, Z => n1813);
   U1118 : BUF_X1 port map( A => n1819, Z => n1824);
   U1119 : BUF_X1 port map( A => n1830, Z => n1835);
   U1120 : BUF_X1 port map( A => n2545, Z => n2550);
   U1121 : BUF_X1 port map( A => n2556, Z => n2561);
   U1122 : BUF_X1 port map( A => n2567, Z => n2572);
   U1123 : BUF_X1 port map( A => n2578, Z => n2583);
   U1124 : BUF_X1 port map( A => n2589, Z => n2594);
   U1125 : BUF_X1 port map( A => n2600, Z => n2605);
   U1126 : BUF_X1 port map( A => n2707, Z => n2712);
   U1127 : BUF_X1 port map( A => n2718, Z => n2723);
   U1128 : BUF_X1 port map( A => n2729, Z => n2734);
   U1129 : BUF_X1 port map( A => n2740, Z => n2745);
   U1130 : BUF_X1 port map( A => n2751, Z => n2756);
   U1131 : BUF_X1 port map( A => n2762, Z => n2767);
   U1132 : BUF_X1 port map( A => n2773, Z => n2778);
   U1133 : BUF_X1 port map( A => n2784, Z => n2789);
   U1134 : BUF_X1 port map( A => n2795, Z => n2800);
   U1135 : BUF_X1 port map( A => n2806, Z => n2811);
   U1136 : BUF_X1 port map( A => n2817, Z => n2822);
   U1137 : BUF_X1 port map( A => n2828, Z => n2833);
   U1138 : BUF_X1 port map( A => n2839, Z => n2844);
   U1139 : BUF_X1 port map( A => n2850, Z => n2855);
   U1140 : BUF_X1 port map( A => n2861, Z => n2866);
   U1141 : BUF_X1 port map( A => n2872, Z => n2877);
   U1142 : BUF_X1 port map( A => n2883, Z => n2888);
   U1143 : BUF_X1 port map( A => n2894, Z => n2900);
   U1144 : BUF_X1 port map( A => n2906, Z => n2911);
   U1145 : BUF_X1 port map( A => n2922, Z => n2927);
   U1146 : BUF_X1 port map( A => n2933, Z => n2938);
   U1147 : BUF_X1 port map( A => n2944, Z => n2949);
   U1148 : BUF_X1 port map( A => n1798, Z => n1803);
   U1149 : BUF_X1 port map( A => n1809, Z => n1814);
   U1150 : BUF_X1 port map( A => n1820, Z => n1825);
   U1151 : BUF_X1 port map( A => n1831, Z => n1836);
   U1152 : BUF_X1 port map( A => n2546, Z => n2551);
   U1153 : BUF_X1 port map( A => n2557, Z => n2562);
   U1154 : BUF_X1 port map( A => n2568, Z => n2573);
   U1155 : BUF_X1 port map( A => n2579, Z => n2584);
   U1156 : BUF_X1 port map( A => n2590, Z => n2595);
   U1157 : BUF_X1 port map( A => n2601, Z => n2606);
   U1158 : BUF_X1 port map( A => n2708, Z => n2713);
   U1159 : BUF_X1 port map( A => n2719, Z => n2724);
   U1160 : BUF_X1 port map( A => n2730, Z => n2735);
   U1161 : BUF_X1 port map( A => n2741, Z => n2746);
   U1162 : BUF_X1 port map( A => n2752, Z => n2757);
   U1163 : BUF_X1 port map( A => n2763, Z => n2768);
   U1164 : BUF_X1 port map( A => n2774, Z => n2779);
   U1165 : BUF_X1 port map( A => n2785, Z => n2790);
   U1166 : BUF_X1 port map( A => n2796, Z => n2801);
   U1167 : BUF_X1 port map( A => n2807, Z => n2812);
   U1168 : BUF_X1 port map( A => n2818, Z => n2823);
   U1169 : BUF_X1 port map( A => n2829, Z => n2834);
   U1170 : BUF_X1 port map( A => n2840, Z => n2845);
   U1171 : BUF_X1 port map( A => n2851, Z => n2856);
   U1172 : BUF_X1 port map( A => n2862, Z => n2867);
   U1173 : BUF_X1 port map( A => n2873, Z => n2878);
   U1174 : BUF_X1 port map( A => n2884, Z => n2889);
   U1175 : BUF_X1 port map( A => n2895, Z => n2901);
   U1176 : BUF_X1 port map( A => n2907, Z => n2912);
   U1177 : BUF_X1 port map( A => n2923, Z => n2928);
   U1178 : BUF_X1 port map( A => n2934, Z => n2939);
   U1179 : BUF_X1 port map( A => n2945, Z => n2950);
   U1180 : BUF_X1 port map( A => n1798, Z => n1804);
   U1181 : BUF_X1 port map( A => n1809, Z => n1815);
   U1182 : BUF_X1 port map( A => n1820, Z => n1826);
   U1183 : BUF_X1 port map( A => n1831, Z => n1837);
   U1184 : BUF_X1 port map( A => n2546, Z => n2552);
   U1185 : BUF_X1 port map( A => n2557, Z => n2563);
   U1186 : BUF_X1 port map( A => n2568, Z => n2574);
   U1187 : BUF_X1 port map( A => n2579, Z => n2585);
   U1188 : BUF_X1 port map( A => n2590, Z => n2596);
   U1189 : BUF_X1 port map( A => n2601, Z => n2607);
   U1190 : BUF_X1 port map( A => n2708, Z => n2714);
   U1191 : BUF_X1 port map( A => n2719, Z => n2725);
   U1192 : BUF_X1 port map( A => n2730, Z => n2736);
   U1193 : BUF_X1 port map( A => n2741, Z => n2747);
   U1194 : BUF_X1 port map( A => n2752, Z => n2758);
   U1195 : BUF_X1 port map( A => n2763, Z => n2769);
   U1196 : BUF_X1 port map( A => n2774, Z => n2780);
   U1197 : BUF_X1 port map( A => n2785, Z => n2791);
   U1198 : BUF_X1 port map( A => n2796, Z => n2802);
   U1199 : BUF_X1 port map( A => n2807, Z => n2813);
   U1200 : BUF_X1 port map( A => n2818, Z => n2824);
   U1201 : BUF_X1 port map( A => n2829, Z => n2835);
   U1202 : BUF_X1 port map( A => n2840, Z => n2846);
   U1203 : BUF_X1 port map( A => n2851, Z => n2857);
   U1204 : BUF_X1 port map( A => n2862, Z => n2868);
   U1205 : BUF_X1 port map( A => n2873, Z => n2879);
   U1206 : BUF_X1 port map( A => n2884, Z => n2890);
   U1207 : BUF_X1 port map( A => n2895, Z => n2902);
   U1208 : BUF_X1 port map( A => n2907, Z => n2913);
   U1209 : BUF_X1 port map( A => n2923, Z => n2929);
   U1210 : BUF_X1 port map( A => n2934, Z => n2940);
   U1211 : BUF_X1 port map( A => n2945, Z => n2951);
   U1212 : BUF_X1 port map( A => n1798, Z => n1805);
   U1213 : BUF_X1 port map( A => n1809, Z => n1816);
   U1214 : BUF_X1 port map( A => n1820, Z => n1827);
   U1215 : BUF_X1 port map( A => n1831, Z => n1838);
   U1216 : BUF_X1 port map( A => n2546, Z => n2553);
   U1217 : BUF_X1 port map( A => n2557, Z => n2564);
   U1218 : BUF_X1 port map( A => n2568, Z => n2575);
   U1219 : BUF_X1 port map( A => n2579, Z => n2586);
   U1220 : BUF_X1 port map( A => n2590, Z => n2597);
   U1221 : BUF_X1 port map( A => n2601, Z => n2704);
   U1222 : BUF_X1 port map( A => n2708, Z => n2715);
   U1223 : BUF_X1 port map( A => n2719, Z => n2726);
   U1224 : BUF_X1 port map( A => n2730, Z => n2737);
   U1225 : BUF_X1 port map( A => n2741, Z => n2748);
   U1226 : BUF_X1 port map( A => n2752, Z => n2759);
   U1227 : BUF_X1 port map( A => n2763, Z => n2770);
   U1228 : BUF_X1 port map( A => n2774, Z => n2781);
   U1229 : BUF_X1 port map( A => n2785, Z => n2792);
   U1230 : BUF_X1 port map( A => n2796, Z => n2803);
   U1231 : BUF_X1 port map( A => n2807, Z => n2814);
   U1232 : BUF_X1 port map( A => n2818, Z => n2825);
   U1233 : BUF_X1 port map( A => n2829, Z => n2836);
   U1234 : BUF_X1 port map( A => n2840, Z => n2847);
   U1235 : BUF_X1 port map( A => n2851, Z => n2858);
   U1236 : BUF_X1 port map( A => n2862, Z => n2869);
   U1237 : BUF_X1 port map( A => n2873, Z => n2880);
   U1238 : BUF_X1 port map( A => n2884, Z => n2891);
   U1239 : BUF_X1 port map( A => n2895, Z => n2903);
   U1240 : BUF_X1 port map( A => n2907, Z => n2914);
   U1241 : BUF_X1 port map( A => n2923, Z => n2930);
   U1242 : BUF_X1 port map( A => n2934, Z => n2941);
   U1243 : BUF_X1 port map( A => n2945, Z => n2952);
   U1244 : BUF_X1 port map( A => n1799, Z => n1806);
   U1245 : BUF_X1 port map( A => n1810, Z => n1817);
   U1246 : BUF_X1 port map( A => n1821, Z => n1828);
   U1247 : BUF_X1 port map( A => n1832, Z => n1839);
   U1248 : BUF_X1 port map( A => n2547, Z => n2554);
   U1249 : BUF_X1 port map( A => n2558, Z => n2565);
   U1250 : BUF_X1 port map( A => n2569, Z => n2576);
   U1251 : BUF_X1 port map( A => n2580, Z => n2587);
   U1252 : BUF_X1 port map( A => n2591, Z => n2598);
   U1253 : BUF_X1 port map( A => n2602, Z => n2705);
   U1254 : BUF_X1 port map( A => n2709, Z => n2716);
   U1255 : BUF_X1 port map( A => n2720, Z => n2727);
   U1256 : BUF_X1 port map( A => n2731, Z => n2738);
   U1257 : BUF_X1 port map( A => n2742, Z => n2749);
   U1258 : BUF_X1 port map( A => n2753, Z => n2760);
   U1259 : BUF_X1 port map( A => n2764, Z => n2771);
   U1260 : BUF_X1 port map( A => n2775, Z => n2782);
   U1261 : BUF_X1 port map( A => n2786, Z => n2793);
   U1262 : BUF_X1 port map( A => n2797, Z => n2804);
   U1263 : BUF_X1 port map( A => n2808, Z => n2815);
   U1264 : BUF_X1 port map( A => n2819, Z => n2826);
   U1265 : BUF_X1 port map( A => n2830, Z => n2837);
   U1266 : BUF_X1 port map( A => n2841, Z => n2848);
   U1267 : BUF_X1 port map( A => n2852, Z => n2859);
   U1268 : BUF_X1 port map( A => n2863, Z => n2870);
   U1269 : BUF_X1 port map( A => n2874, Z => n2881);
   U1270 : BUF_X1 port map( A => n2885, Z => n2892);
   U1271 : BUF_X1 port map( A => n2896, Z => n2904);
   U1272 : BUF_X1 port map( A => n2908, Z => n2915);
   U1273 : BUF_X1 port map( A => n2924, Z => n2931);
   U1274 : BUF_X1 port map( A => n2935, Z => n2942);
   U1275 : BUF_X1 port map( A => n2946, Z => n2953);
   U1276 : BUF_X1 port map( A => n1799, Z => n1807);
   U1277 : BUF_X1 port map( A => n1810, Z => n1818);
   U1278 : BUF_X1 port map( A => n1821, Z => n1829);
   U1279 : BUF_X1 port map( A => n1832, Z => n2544);
   U1280 : BUF_X1 port map( A => n2547, Z => n2555);
   U1281 : BUF_X1 port map( A => n2558, Z => n2566);
   U1282 : BUF_X1 port map( A => n2569, Z => n2577);
   U1283 : BUF_X1 port map( A => n2580, Z => n2588);
   U1284 : BUF_X1 port map( A => n2591, Z => n2599);
   U1285 : BUF_X1 port map( A => n2602, Z => n2706);
   U1286 : BUF_X1 port map( A => n2709, Z => n2717);
   U1287 : BUF_X1 port map( A => n2720, Z => n2728);
   U1288 : BUF_X1 port map( A => n2731, Z => n2739);
   U1289 : BUF_X1 port map( A => n2742, Z => n2750);
   U1290 : BUF_X1 port map( A => n2753, Z => n2761);
   U1291 : BUF_X1 port map( A => n2764, Z => n2772);
   U1292 : BUF_X1 port map( A => n2775, Z => n2783);
   U1293 : BUF_X1 port map( A => n2786, Z => n2794);
   U1294 : BUF_X1 port map( A => n2797, Z => n2805);
   U1295 : BUF_X1 port map( A => n2808, Z => n2816);
   U1296 : BUF_X1 port map( A => n2819, Z => n2827);
   U1297 : BUF_X1 port map( A => n2830, Z => n2838);
   U1298 : BUF_X1 port map( A => n2841, Z => n2849);
   U1299 : BUF_X1 port map( A => n2852, Z => n2860);
   U1300 : BUF_X1 port map( A => n2863, Z => n2871);
   U1301 : BUF_X1 port map( A => n2874, Z => n2882);
   U1302 : BUF_X1 port map( A => n2885, Z => n2893);
   U1303 : BUF_X1 port map( A => n2896, Z => n2905);
   U1304 : BUF_X1 port map( A => n2908, Z => n2917);
   U1305 : BUF_X1 port map( A => n2924, Z => n2932);
   U1306 : BUF_X1 port map( A => n2935, Z => n2943);
   U1307 : BUF_X1 port map( A => n2946, Z => n2954);
   U1308 : NAND2_X1 port map( A1 => n6247, A2 => n6313, ZN => n4994);
   U1309 : NAND2_X1 port map( A1 => n4804, A2 => n4870, ZN => n3551);
   U1310 : AND2_X1 port map( A1 => n6252, A2 => n6254, ZN => n6248);
   U1311 : AND2_X1 port map( A1 => n6252, A2 => n6253, ZN => n6246);
   U1312 : AND2_X1 port map( A1 => n4809, A2 => n4811, ZN => n4805);
   U1313 : AND2_X1 port map( A1 => n4809, A2 => n4810, ZN => n4803);
   U1314 : AND2_X1 port map( A1 => n6254, A2 => n6297, ZN => n6298);
   U1315 : AND2_X1 port map( A1 => n4811, A2 => n4854, ZN => n4855);
   U1316 : NAND2_X1 port map( A1 => n6297, A2 => n6287, ZN => n4987);
   U1317 : NAND2_X1 port map( A1 => n4854, A2 => n4844, ZN => n3544);
   U1318 : NAND2_X1 port map( A1 => n6283, A2 => n6284, ZN => n4934);
   U1319 : NAND2_X1 port map( A1 => n6283, A2 => n6285, ZN => n4933);
   U1320 : NAND2_X1 port map( A1 => n6283, A2 => n6261, ZN => n4965);
   U1321 : NAND2_X1 port map( A1 => n6283, A2 => n6260, ZN => n4963);
   U1322 : NAND2_X1 port map( A1 => n4840, A2 => n4841, ZN => n3491);
   U1323 : NAND2_X1 port map( A1 => n4840, A2 => n4842, ZN => n3490);
   U1324 : NAND2_X1 port map( A1 => n4840, A2 => n4818, ZN => n3522);
   U1325 : NAND2_X1 port map( A1 => n4840, A2 => n4817, ZN => n3520);
   U1326 : NAND2_X1 port map( A1 => n6255, A2 => n3374, ZN => n4985);
   U1327 : NAND2_X1 port map( A1 => n6257, A2 => n3374, ZN => n4986);
   U1328 : NAND2_X1 port map( A1 => n6256, A2 => n3374, ZN => n4990);
   U1329 : NAND2_X1 port map( A1 => n6262, A2 => n3374, ZN => n4988);
   U1330 : NAND2_X1 port map( A1 => n6263, A2 => n3374, ZN => n4989);
   U1331 : NAND2_X1 port map( A1 => n6260, A2 => n3374, ZN => n4996);
   U1332 : NAND2_X1 port map( A1 => n4812, A2 => n3384, ZN => n3542);
   U1333 : NAND2_X1 port map( A1 => n4814, A2 => n3384, ZN => n3543);
   U1334 : NAND2_X1 port map( A1 => n4813, A2 => n3384, ZN => n3547);
   U1335 : NAND2_X1 port map( A1 => n4819, A2 => n3384, ZN => n3545);
   U1336 : NAND2_X1 port map( A1 => n4820, A2 => n3384, ZN => n3546);
   U1337 : NAND2_X1 port map( A1 => n4817, A2 => n3384, ZN => n3553);
   U1338 : NAND2_X1 port map( A1 => n6252, A2 => n6255, ZN => n4897);
   U1339 : NAND2_X1 port map( A1 => n6252, A2 => n6257, ZN => n4895);
   U1340 : NAND2_X1 port map( A1 => n6252, A2 => n6256, ZN => n4896);
   U1341 : NAND2_X1 port map( A1 => n6252, A2 => n6259, ZN => n4903);
   U1342 : NAND2_X1 port map( A1 => n6252, A2 => n6261, ZN => n4901);
   U1343 : NAND2_X1 port map( A1 => n6252, A2 => n6260, ZN => n4902);
   U1344 : NAND2_X1 port map( A1 => n4809, A2 => n4812, ZN => n3454);
   U1345 : NAND2_X1 port map( A1 => n4809, A2 => n4814, ZN => n3452);
   U1346 : NAND2_X1 port map( A1 => n4809, A2 => n4813, ZN => n3453);
   U1347 : NAND2_X1 port map( A1 => n4809, A2 => n4816, ZN => n3460);
   U1348 : NAND2_X1 port map( A1 => n4809, A2 => n4818, ZN => n3458);
   U1349 : NAND2_X1 port map( A1 => n4809, A2 => n4817, ZN => n3459);
   U1350 : NAND2_X1 port map( A1 => n6248, A2 => n6251, ZN => n4892);
   U1351 : NAND2_X1 port map( A1 => n6246, A2 => n6251, ZN => n4893);
   U1352 : NAND2_X1 port map( A1 => n6267, A2 => n6251, ZN => n4918);
   U1353 : NAND2_X1 port map( A1 => n6268, A2 => n6251, ZN => n4919);
   U1354 : NAND2_X1 port map( A1 => n6298, A2 => n6251, ZN => n4983);
   U1355 : NAND2_X1 port map( A1 => n4805, A2 => n4808, ZN => n3449);
   U1356 : NAND2_X1 port map( A1 => n4803, A2 => n4808, ZN => n3450);
   U1357 : NAND2_X1 port map( A1 => n4824, A2 => n4808, ZN => n3475);
   U1358 : NAND2_X1 port map( A1 => n4825, A2 => n4808, ZN => n3476);
   U1359 : NAND2_X1 port map( A1 => n4855, A2 => n4808, ZN => n3540);
   U1360 : NAND2_X1 port map( A1 => n6248, A2 => n6250, ZN => n4890);
   U1361 : NAND2_X1 port map( A1 => n6246, A2 => n6250, ZN => n4894);
   U1362 : NAND2_X1 port map( A1 => n6281, A2 => n6250, ZN => n4932);
   U1363 : NAND2_X1 port map( A1 => n6298, A2 => n6250, ZN => n4984);
   U1364 : NAND2_X1 port map( A1 => n4805, A2 => n4807, ZN => n3447);
   U1365 : NAND2_X1 port map( A1 => n4803, A2 => n4807, ZN => n3451);
   U1366 : NAND2_X1 port map( A1 => n4838, A2 => n4807, ZN => n3489);
   U1367 : NAND2_X1 port map( A1 => n4855, A2 => n4807, ZN => n3541);
   U1368 : AND2_X1 port map( A1 => n6283, A2 => n6254, ZN => n6281);
   U1369 : AND2_X1 port map( A1 => n4840, A2 => n4811, ZN => n4838);
   U1370 : NAND2_X1 port map( A1 => n6286, A2 => n6297, ZN => n4958);
   U1371 : NAND2_X1 port map( A1 => n6285, A2 => n6297, ZN => n4982);
   U1372 : NAND2_X1 port map( A1 => n6284, A2 => n6297, ZN => n4981);
   U1373 : NAND2_X1 port map( A1 => n4843, A2 => n4854, ZN => n3515);
   U1374 : NAND2_X1 port map( A1 => n4842, A2 => n4854, ZN => n3539);
   U1375 : NAND2_X1 port map( A1 => n4841, A2 => n4854, ZN => n3538);
   U1376 : BUF_X1 port map( A => RESET, Z => n2955);
   U1377 : NAND2_X1 port map( A1 => n6279, A2 => n6260, ZN => n4926);
   U1378 : NAND2_X1 port map( A1 => n4836, A2 => n4817, ZN => n3483);
   U1379 : NAND2_X1 port map( A1 => n6279, A2 => n6261, ZN => n4928);
   U1380 : NAND2_X1 port map( A1 => n4836, A2 => n4818, ZN => n3485);
   U1381 : NAND2_X1 port map( A1 => n6279, A2 => n6256, ZN => n4921);
   U1382 : NAND2_X1 port map( A1 => n4836, A2 => n4813, ZN => n3478);
   U1383 : NAND2_X1 port map( A1 => n6279, A2 => n6255, ZN => n4922);
   U1384 : NAND2_X1 port map( A1 => n6279, A2 => n6257, ZN => n4920);
   U1385 : NAND2_X1 port map( A1 => n4836, A2 => n4812, ZN => n3479);
   U1386 : NAND2_X1 port map( A1 => n4836, A2 => n4814, ZN => n3477);
   U1387 : NAND2_X1 port map( A1 => n6279, A2 => n6259, ZN => n4924);
   U1388 : NAND2_X1 port map( A1 => n4836, A2 => n4816, ZN => n3481);
   U1389 : NAND2_X1 port map( A1 => n6279, A2 => n6262, ZN => n4925);
   U1390 : NAND2_X1 port map( A1 => n4836, A2 => n4819, ZN => n3482);
   U1391 : NAND2_X1 port map( A1 => n6279, A2 => n6263, ZN => n4923);
   U1392 : NAND2_X1 port map( A1 => n4836, A2 => n4820, ZN => n3480);
   U1393 : AND2_X1 port map( A1 => n6249, A2 => n6312, ZN => n5002);
   U1394 : AND2_X1 port map( A1 => n6249, A2 => n6313, ZN => n5000);
   U1395 : AND2_X1 port map( A1 => n4806, A2 => n4869, ZN => n3559);
   U1396 : AND2_X1 port map( A1 => n4806, A2 => n4870, ZN => n3557);
   U1397 : AND2_X1 port map( A1 => n6296, A2 => n6254, ZN => n6300);
   U1398 : AND2_X1 port map( A1 => n4853, A2 => n4811, ZN => n4857);
   U1399 : AND2_X1 port map( A1 => n6316, A2 => n3381, ZN => n6312);
   U1400 : AND2_X1 port map( A1 => n4873, A2 => n3389, ZN => n4869);
   U1401 : AND2_X1 port map( A1 => n6253, A2 => n6249, ZN => n6284);
   U1402 : AND2_X1 port map( A1 => n4810, A2 => n4806, ZN => n4841);
   U1403 : AND2_X1 port map( A1 => n6268, A2 => n6249, ZN => n4904);
   U1404 : AND2_X1 port map( A1 => n6267, A2 => n6249, ZN => n4908);
   U1405 : AND2_X1 port map( A1 => n6281, A2 => n6249, ZN => n4929);
   U1406 : AND2_X1 port map( A1 => n6300, A2 => n6249, ZN => n4971);
   U1407 : AND2_X1 port map( A1 => n4825, A2 => n4806, ZN => n3461);
   U1408 : AND2_X1 port map( A1 => n4824, A2 => n4806, ZN => n3465);
   U1409 : AND2_X1 port map( A1 => n4838, A2 => n4806, ZN => n3486);
   U1410 : AND2_X1 port map( A1 => n4857, A2 => n4806, ZN => n3528);
   U1411 : AND2_X1 port map( A1 => n6253, A2 => n6251, ZN => n6287);
   U1412 : AND2_X1 port map( A1 => n4810, A2 => n4808, ZN => n4844);
   U1413 : AND2_X1 port map( A1 => n6296, A2 => n6285, ZN => n4968);
   U1414 : AND2_X1 port map( A1 => n6296, A2 => n6284, ZN => n4970);
   U1415 : AND2_X1 port map( A1 => n6296, A2 => n6286, ZN => n4969);
   U1416 : AND2_X1 port map( A1 => n4853, A2 => n4842, ZN => n3525);
   U1417 : AND2_X1 port map( A1 => n4853, A2 => n4841, ZN => n3527);
   U1418 : AND2_X1 port map( A1 => n4853, A2 => n4843, ZN => n3526);
   U1419 : AND2_X1 port map( A1 => n6251, A2 => n6312, ZN => n4998);
   U1420 : AND2_X1 port map( A1 => n4808, A2 => n4869, ZN => n3555);
   U1421 : AND2_X1 port map( A1 => n6283, A2 => n6262, ZN => n4936);
   U1422 : AND2_X1 port map( A1 => n6283, A2 => n6256, ZN => n4937);
   U1423 : AND2_X1 port map( A1 => n6283, A2 => n6257, ZN => n4935);
   U1424 : AND2_X1 port map( A1 => n6283, A2 => n6255, ZN => n4939);
   U1425 : AND2_X1 port map( A1 => n6283, A2 => n6287, ZN => n4940);
   U1426 : AND2_X1 port map( A1 => n6283, A2 => n6286, ZN => n4930);
   U1427 : AND2_X1 port map( A1 => n6283, A2 => n6259, ZN => n4960);
   U1428 : AND2_X1 port map( A1 => n6283, A2 => n6263, ZN => n4961);
   U1429 : AND2_X1 port map( A1 => n4840, A2 => n4819, ZN => n3493);
   U1430 : AND2_X1 port map( A1 => n4840, A2 => n4813, ZN => n3494);
   U1431 : AND2_X1 port map( A1 => n4840, A2 => n4814, ZN => n3492);
   U1432 : AND2_X1 port map( A1 => n4840, A2 => n4812, ZN => n3496);
   U1433 : AND2_X1 port map( A1 => n4840, A2 => n4844, ZN => n3497);
   U1434 : AND2_X1 port map( A1 => n4840, A2 => n4843, ZN => n3487);
   U1435 : AND2_X1 port map( A1 => n4840, A2 => n4816, ZN => n3517);
   U1436 : AND2_X1 port map( A1 => n4840, A2 => n4820, ZN => n3518);
   U1437 : AND2_X1 port map( A1 => n6250, A2 => n6312, ZN => n4997);
   U1438 : AND2_X1 port map( A1 => n6250, A2 => n6313, ZN => n5001);
   U1439 : AND2_X1 port map( A1 => n4807, A2 => n4869, ZN => n3554);
   U1440 : AND2_X1 port map( A1 => n4807, A2 => n4870, ZN => n3558);
   U1441 : AND2_X1 port map( A1 => n6267, A2 => n6247, ZN => n4907);
   U1442 : AND2_X1 port map( A1 => n4824, A2 => n4804, ZN => n3464);
   U1443 : AND2_X1 port map( A1 => n6252, A2 => n6263, ZN => n4898);
   U1444 : AND2_X1 port map( A1 => n6252, A2 => n6262, ZN => n4899);
   U1445 : AND2_X1 port map( A1 => n4809, A2 => n4820, ZN => n3455);
   U1446 : AND2_X1 port map( A1 => n4809, A2 => n4819, ZN => n3456);
   U1447 : AND2_X1 port map( A1 => n6281, A2 => n6251, ZN => n4938);
   U1448 : AND2_X1 port map( A1 => n6300, A2 => n6251, ZN => n4967);
   U1449 : AND2_X1 port map( A1 => n6313, A2 => n6251, ZN => n4999);
   U1450 : AND2_X1 port map( A1 => n4838, A2 => n4808, ZN => n3495);
   U1451 : AND2_X1 port map( A1 => n4857, A2 => n4808, ZN => n3524);
   U1452 : AND2_X1 port map( A1 => n4870, A2 => n4808, ZN => n3556);
   U1453 : AND2_X1 port map( A1 => n6253, A2 => n6250, ZN => n6285);
   U1454 : AND2_X1 port map( A1 => n4810, A2 => n4807, ZN => n4842);
   U1455 : AND2_X1 port map( A1 => n6268, A2 => n6250, ZN => n4905);
   U1456 : AND2_X1 port map( A1 => n6267, A2 => n6250, ZN => n4906);
   U1457 : AND2_X1 port map( A1 => n6300, A2 => n6250, ZN => n4966);
   U1458 : AND2_X1 port map( A1 => n4825, A2 => n4807, ZN => n3462);
   U1459 : AND2_X1 port map( A1 => n4824, A2 => n4807, ZN => n3463);
   U1460 : AND2_X1 port map( A1 => n4857, A2 => n4807, ZN => n3523);
   U1461 : AND2_X1 port map( A1 => n6277, A2 => n3381, ZN => n6268);
   U1462 : AND2_X1 port map( A1 => n4834, A2 => n3389, ZN => n4825);
   U1463 : AND2_X1 port map( A1 => n6261, A2 => n3374, ZN => n4991);
   U1464 : AND2_X1 port map( A1 => n6259, A2 => n3374, ZN => n4992);
   U1465 : AND2_X1 port map( A1 => n4818, A2 => n3384, ZN => n3548);
   U1466 : AND2_X1 port map( A1 => n4816, A2 => n3384, ZN => n3549);
   U1467 : AND2_X1 port map( A1 => n6253, A2 => n6247, ZN => n6286);
   U1468 : AND2_X1 port map( A1 => n4810, A2 => n4804, ZN => n4843);
   U1469 : INV_X1 port map( A => n3419, ZN => n3392);
   U1470 : NAND4_X1 port map( A1 => n3106, A2 => n3108, A3 => n3368, A4 => 
                           n3365, ZN => n3382);
   U1471 : NOR2_X1 port map( A1 => n3376, A2 => n6266, ZN => n6297);
   U1472 : NOR2_X1 port map( A1 => n3385, A2 => n4823, ZN => n4854);
   U1473 : NOR2_X1 port map( A1 => n3405, A2 => n3406, ZN => n3358);
   U1474 : NOR2_X1 port map( A1 => n3373, A2 => n3406, ZN => n3353);
   U1475 : NOR2_X1 port map( A1 => n3372, A2 => n3405, ZN => n3348);
   U1476 : NOR2_X1 port map( A1 => n3377, A2 => n3359, ZN => n3364);
   U1477 : NOR2_X1 port map( A1 => n3370, A2 => n3359, ZN => n3342);
   U1478 : NOR2_X1 port map( A1 => n3369, A2 => n3377, ZN => n3400);
   U1479 : INV_X1 port map( A => N8415, ZN => n10918);
   U1480 : INV_X1 port map( A => N8559, ZN => n10919);
   U1481 : INV_X1 port map( A => N2151, ZN => n3391);
   U1482 : AND3_X1 port map( A1 => n6264, A2 => n6265, A3 => n6266, ZN => n6252
                           );
   U1483 : AND3_X1 port map( A1 => n4821, A2 => n4822, A3 => n4823, ZN => n4809
                           );
   U1484 : INV_X1 port map( A => n6266, ZN => n3374);
   U1485 : INV_X1 port map( A => n4823, ZN => n3384);
   U1486 : NOR2_X1 port map( A1 => n6278, A2 => n6280, ZN => n6309);
   U1487 : NOR2_X1 port map( A1 => n4835, A2 => n4837, ZN => n4866);
   U1488 : NOR2_X1 port map( A1 => n3381, A2 => n6280, ZN => n6310);
   U1489 : NOR2_X1 port map( A1 => n3389, A2 => n4837, ZN => n4867);
   U1490 : INV_X1 port map( A => n3109, ZN => n3368);
   U1491 : INV_X1 port map( A => n3108, ZN => n3366);
   U1492 : INV_X1 port map( A => n3107, ZN => n3365);
   U1493 : AND2_X1 port map( A1 => n6264, A2 => n3376, ZN => n6279);
   U1494 : AND2_X1 port map( A1 => n4821, A2 => n3385, ZN => n4836);
   U1495 : INV_X1 port map( A => n6265, ZN => n3376);
   U1496 : INV_X1 port map( A => n4822, ZN => n3385);
   U1497 : INV_X1 port map( A => n6314, ZN => n3379);
   U1498 : INV_X1 port map( A => n4871, ZN => n3388);
   U1499 : NOR2_X1 port map( A1 => n6265, A2 => n6266, ZN => n6316);
   U1500 : NOR2_X1 port map( A1 => n4822, A2 => n4823, ZN => n4873);
   U1501 : INV_X1 port map( A => n6315, ZN => n3378);
   U1502 : INV_X1 port map( A => n4872, ZN => n3387);
   U1503 : INV_X1 port map( A => n6278, ZN => n3381);
   U1504 : INV_X1 port map( A => n4835, ZN => n3389);
   U1505 : AND2_X1 port map( A1 => n6280, A2 => n3381, ZN => n6253);
   U1506 : AND2_X1 port map( A1 => n4837, A2 => n3389, ZN => n4810);
   U1507 : AND2_X1 port map( A1 => n6278, A2 => n6316, ZN => n6313);
   U1508 : AND2_X1 port map( A1 => n4835, A2 => n4873, ZN => n4870);
   U1509 : BUF_X1 port map( A => N8702, Z => n1795);
   U1510 : BUF_X1 port map( A => N8735, Z => n1792);
   U1511 : BUF_X1 port map( A => N8702, Z => n1794);
   U1512 : BUF_X1 port map( A => N8735, Z => n1791);
   U1513 : AND2_X1 port map( A1 => n6277, A2 => n6278, ZN => n6267);
   U1514 : AND2_X1 port map( A1 => n4834, A2 => n4835, ZN => n4824);
   U1515 : BUF_X1 port map( A => N8702, Z => n1796);
   U1516 : BUF_X1 port map( A => N8735, Z => n1793);
   U1517 : AND2_X1 port map( A1 => n6280, A2 => n6278, ZN => n6254);
   U1518 : AND2_X1 port map( A1 => n4837, A2 => n4835, ZN => n4811);
   U1519 : INV_X1 port map( A => n3405, ZN => n3373);
   U1520 : INV_X1 port map( A => n3377, ZN => n3370);
   U1521 : INV_X1 port map( A => n3406, ZN => n3372);
   U1522 : INV_X1 port map( A => n3359, ZN => n3369);
   U1523 : AND3_X1 port map( A1 => n6279, A2 => n6280, A3 => n6266, ZN => n6277
                           );
   U1524 : AND3_X1 port map( A1 => n4836, A2 => n4837, A3 => n4823, ZN => n4834
                           );
   U1525 : NOR2_X1 port map( A1 => n3265, A2 => n6233, ZN => N8703);
   U1526 : NOR4_X1 port map( A1 => n6234, A2 => n6235, A3 => n6236, A4 => n6237
                           , ZN => n6233);
   U1527 : NAND4_X1 port map( A1 => n6301, A2 => n6302, A3 => n6303, A4 => 
                           n6304, ZN => n6234);
   U1528 : NAND4_X1 port map( A1 => n6288, A2 => n6289, A3 => n6290, A4 => 
                           n6291, ZN => n6235);
   U1529 : NOR2_X1 port map( A1 => n3276, A2 => n4790, ZN => N8736);
   U1530 : NOR4_X1 port map( A1 => n4791, A2 => n4792, A3 => n4793, A4 => n4794
                           , ZN => n4790);
   U1531 : NAND4_X1 port map( A1 => n4858, A2 => n4859, A3 => n4860, A4 => 
                           n4861, ZN => n4791);
   U1532 : NAND4_X1 port map( A1 => n4845, A2 => n4846, A3 => n4847, A4 => 
                           n4848, ZN => n4792);
   U1533 : NOR2_X1 port map( A1 => n3265, A2 => n6192, ZN => N8704);
   U1534 : NOR4_X1 port map( A1 => n6193, A2 => n6194, A3 => n6195, A4 => n6196
                           , ZN => n6192);
   U1535 : NAND4_X1 port map( A1 => n6224, A2 => n6225, A3 => n6226, A4 => 
                           n6227, ZN => n6193);
   U1536 : NAND4_X1 port map( A1 => n6215, A2 => n6216, A3 => n6217, A4 => 
                           n6218, ZN => n6194);
   U1537 : NOR2_X1 port map( A1 => n3276, A2 => n4749, ZN => N8737);
   U1538 : NOR4_X1 port map( A1 => n4750, A2 => n4751, A3 => n4752, A4 => n4753
                           , ZN => n4749);
   U1539 : NAND4_X1 port map( A1 => n4781, A2 => n4782, A3 => n4783, A4 => 
                           n4784, ZN => n4750);
   U1540 : NAND4_X1 port map( A1 => n4772, A2 => n4773, A3 => n4774, A4 => 
                           n4775, ZN => n4751);
   U1541 : NOR2_X1 port map( A1 => n3265, A2 => n6151, ZN => N8705);
   U1542 : NOR4_X1 port map( A1 => n6152, A2 => n6153, A3 => n6154, A4 => n6155
                           , ZN => n6151);
   U1543 : NAND4_X1 port map( A1 => n6183, A2 => n6184, A3 => n6185, A4 => 
                           n6186, ZN => n6152);
   U1544 : NAND4_X1 port map( A1 => n6174, A2 => n6175, A3 => n6176, A4 => 
                           n6177, ZN => n6153);
   U1545 : NOR2_X1 port map( A1 => n3276, A2 => n4708, ZN => N8738);
   U1546 : NOR4_X1 port map( A1 => n4709, A2 => n4710, A3 => n4711, A4 => n4712
                           , ZN => n4708);
   U1547 : NAND4_X1 port map( A1 => n4740, A2 => n4741, A3 => n4742, A4 => 
                           n4743, ZN => n4709);
   U1548 : NAND4_X1 port map( A1 => n4731, A2 => n4732, A3 => n4733, A4 => 
                           n4734, ZN => n4710);
   U1549 : NOR2_X1 port map( A1 => n3265, A2 => n6110, ZN => N8706);
   U1550 : NOR4_X1 port map( A1 => n6111, A2 => n6112, A3 => n6113, A4 => n6114
                           , ZN => n6110);
   U1551 : NAND4_X1 port map( A1 => n6142, A2 => n6143, A3 => n6144, A4 => 
                           n6145, ZN => n6111);
   U1552 : NAND4_X1 port map( A1 => n6133, A2 => n6134, A3 => n6135, A4 => 
                           n6136, ZN => n6112);
   U1553 : NOR2_X1 port map( A1 => n3277, A2 => n4667, ZN => N8739);
   U1554 : NOR4_X1 port map( A1 => n4668, A2 => n4669, A3 => n4670, A4 => n4671
                           , ZN => n4667);
   U1555 : NAND4_X1 port map( A1 => n4699, A2 => n4700, A3 => n4701, A4 => 
                           n4702, ZN => n4668);
   U1556 : NAND4_X1 port map( A1 => n4690, A2 => n4691, A3 => n4692, A4 => 
                           n4693, ZN => n4669);
   U1557 : NOR2_X1 port map( A1 => n3266, A2 => n6069, ZN => N8707);
   U1558 : NOR4_X1 port map( A1 => n6070, A2 => n6071, A3 => n6072, A4 => n6073
                           , ZN => n6069);
   U1559 : NAND4_X1 port map( A1 => n6101, A2 => n6102, A3 => n6103, A4 => 
                           n6104, ZN => n6070);
   U1560 : NAND4_X1 port map( A1 => n6092, A2 => n6093, A3 => n6094, A4 => 
                           n6095, ZN => n6071);
   U1561 : NOR2_X1 port map( A1 => n3277, A2 => n4626, ZN => N8740);
   U1562 : NOR4_X1 port map( A1 => n4627, A2 => n4628, A3 => n4629, A4 => n4630
                           , ZN => n4626);
   U1563 : NAND4_X1 port map( A1 => n4658, A2 => n4659, A3 => n4660, A4 => 
                           n4661, ZN => n4627);
   U1564 : NAND4_X1 port map( A1 => n4649, A2 => n4650, A3 => n4651, A4 => 
                           n4652, ZN => n4628);
   U1565 : NOR2_X1 port map( A1 => n3266, A2 => n6028, ZN => N8708);
   U1566 : NOR4_X1 port map( A1 => n6029, A2 => n6030, A3 => n6031, A4 => n6032
                           , ZN => n6028);
   U1567 : NAND4_X1 port map( A1 => n6060, A2 => n6061, A3 => n6062, A4 => 
                           n6063, ZN => n6029);
   U1568 : NAND4_X1 port map( A1 => n6051, A2 => n6052, A3 => n6053, A4 => 
                           n6054, ZN => n6030);
   U1569 : NOR2_X1 port map( A1 => n3277, A2 => n4585, ZN => N8741);
   U1570 : NOR4_X1 port map( A1 => n4586, A2 => n4587, A3 => n4588, A4 => n4589
                           , ZN => n4585);
   U1571 : NAND4_X1 port map( A1 => n4617, A2 => n4618, A3 => n4619, A4 => 
                           n4620, ZN => n4586);
   U1572 : NAND4_X1 port map( A1 => n4608, A2 => n4609, A3 => n4610, A4 => 
                           n4611, ZN => n4587);
   U1573 : NOR2_X1 port map( A1 => n3266, A2 => n5987, ZN => N8709);
   U1574 : NOR4_X1 port map( A1 => n5988, A2 => n5989, A3 => n5990, A4 => n5991
                           , ZN => n5987);
   U1575 : NAND4_X1 port map( A1 => n6019, A2 => n6020, A3 => n6021, A4 => 
                           n6022, ZN => n5988);
   U1576 : NAND4_X1 port map( A1 => n6010, A2 => n6011, A3 => n6012, A4 => 
                           n6013, ZN => n5989);
   U1577 : NOR2_X1 port map( A1 => n3277, A2 => n4544, ZN => N8742);
   U1578 : NOR4_X1 port map( A1 => n4545, A2 => n4546, A3 => n4547, A4 => n4548
                           , ZN => n4544);
   U1579 : NAND4_X1 port map( A1 => n4576, A2 => n4577, A3 => n4578, A4 => 
                           n4579, ZN => n4545);
   U1580 : NAND4_X1 port map( A1 => n4567, A2 => n4568, A3 => n4569, A4 => 
                           n4570, ZN => n4546);
   U1581 : NOR2_X1 port map( A1 => n3266, A2 => n5946, ZN => N8710);
   U1582 : NOR4_X1 port map( A1 => n5947, A2 => n5948, A3 => n5949, A4 => n5950
                           , ZN => n5946);
   U1583 : NAND4_X1 port map( A1 => n5978, A2 => n5979, A3 => n5980, A4 => 
                           n5981, ZN => n5947);
   U1584 : NAND4_X1 port map( A1 => n5969, A2 => n5970, A3 => n5971, A4 => 
                           n5972, ZN => n5948);
   U1585 : NOR2_X1 port map( A1 => n3278, A2 => n4503, ZN => N8743);
   U1586 : NOR4_X1 port map( A1 => n4504, A2 => n4505, A3 => n4506, A4 => n4507
                           , ZN => n4503);
   U1587 : NAND4_X1 port map( A1 => n4535, A2 => n4536, A3 => n4537, A4 => 
                           n4538, ZN => n4504);
   U1588 : NAND4_X1 port map( A1 => n4526, A2 => n4527, A3 => n4528, A4 => 
                           n4529, ZN => n4505);
   U1589 : NOR2_X1 port map( A1 => n3268, A2 => n5905, ZN => N8711);
   U1590 : NOR4_X1 port map( A1 => n5906, A2 => n5907, A3 => n5908, A4 => n5909
                           , ZN => n5905);
   U1591 : NAND4_X1 port map( A1 => n5937, A2 => n5938, A3 => n5939, A4 => 
                           n5940, ZN => n5906);
   U1592 : NAND4_X1 port map( A1 => n5928, A2 => n5929, A3 => n5930, A4 => 
                           n5931, ZN => n5907);
   U1593 : NOR2_X1 port map( A1 => n3278, A2 => n4462, ZN => N8744);
   U1594 : NOR4_X1 port map( A1 => n4463, A2 => n4464, A3 => n4465, A4 => n4466
                           , ZN => n4462);
   U1595 : NAND4_X1 port map( A1 => n4494, A2 => n4495, A3 => n4496, A4 => 
                           n4497, ZN => n4463);
   U1596 : NAND4_X1 port map( A1 => n4485, A2 => n4486, A3 => n4487, A4 => 
                           n4488, ZN => n4464);
   U1597 : NOR2_X1 port map( A1 => n3268, A2 => n5864, ZN => N8712);
   U1598 : NOR4_X1 port map( A1 => n5865, A2 => n5866, A3 => n5867, A4 => n5868
                           , ZN => n5864);
   U1599 : NAND4_X1 port map( A1 => n5896, A2 => n5897, A3 => n5898, A4 => 
                           n5899, ZN => n5865);
   U1600 : NAND4_X1 port map( A1 => n5887, A2 => n5888, A3 => n5889, A4 => 
                           n5890, ZN => n5866);
   U1601 : NOR2_X1 port map( A1 => n3278, A2 => n4421, ZN => N8745);
   U1602 : NOR4_X1 port map( A1 => n4422, A2 => n4423, A3 => n4424, A4 => n4425
                           , ZN => n4421);
   U1603 : NAND4_X1 port map( A1 => n4453, A2 => n4454, A3 => n4455, A4 => 
                           n4456, ZN => n4422);
   U1604 : NAND4_X1 port map( A1 => n4444, A2 => n4445, A3 => n4446, A4 => 
                           n4447, ZN => n4423);
   U1605 : NOR2_X1 port map( A1 => n3268, A2 => n5823, ZN => N8713);
   U1606 : NOR4_X1 port map( A1 => n5824, A2 => n5825, A3 => n5826, A4 => n5827
                           , ZN => n5823);
   U1607 : NAND4_X1 port map( A1 => n5855, A2 => n5856, A3 => n5857, A4 => 
                           n5858, ZN => n5824);
   U1608 : NAND4_X1 port map( A1 => n5846, A2 => n5847, A3 => n5848, A4 => 
                           n5849, ZN => n5825);
   U1609 : NOR2_X1 port map( A1 => n3278, A2 => n4380, ZN => N8746);
   U1610 : NOR4_X1 port map( A1 => n4381, A2 => n4382, A3 => n4383, A4 => n4384
                           , ZN => n4380);
   U1611 : NAND4_X1 port map( A1 => n4412, A2 => n4413, A3 => n4414, A4 => 
                           n4415, ZN => n4381);
   U1612 : NAND4_X1 port map( A1 => n4403, A2 => n4404, A3 => n4405, A4 => 
                           n4406, ZN => n4382);
   U1613 : NOR2_X1 port map( A1 => n3268, A2 => n5782, ZN => N8714);
   U1614 : NOR4_X1 port map( A1 => n5783, A2 => n5784, A3 => n5785, A4 => n5786
                           , ZN => n5782);
   U1615 : NAND4_X1 port map( A1 => n5814, A2 => n5815, A3 => n5816, A4 => 
                           n5817, ZN => n5783);
   U1616 : NAND4_X1 port map( A1 => n5805, A2 => n5806, A3 => n5807, A4 => 
                           n5808, ZN => n5784);
   U1617 : NOR2_X1 port map( A1 => n3280, A2 => n4339, ZN => N8747);
   U1618 : NOR4_X1 port map( A1 => n4340, A2 => n4341, A3 => n4342, A4 => n4343
                           , ZN => n4339);
   U1619 : NAND4_X1 port map( A1 => n4371, A2 => n4372, A3 => n4373, A4 => 
                           n4374, ZN => n4340);
   U1620 : NAND4_X1 port map( A1 => n4362, A2 => n4363, A3 => n4364, A4 => 
                           n4365, ZN => n4341);
   U1621 : NOR2_X1 port map( A1 => n3269, A2 => n5741, ZN => N8715);
   U1622 : NOR4_X1 port map( A1 => n5742, A2 => n5743, A3 => n5744, A4 => n5745
                           , ZN => n5741);
   U1623 : NAND4_X1 port map( A1 => n5773, A2 => n5774, A3 => n5775, A4 => 
                           n5776, ZN => n5742);
   U1624 : NAND4_X1 port map( A1 => n5764, A2 => n5765, A3 => n5766, A4 => 
                           n5767, ZN => n5743);
   U1625 : NOR2_X1 port map( A1 => n3280, A2 => n4298, ZN => N8748);
   U1626 : NOR4_X1 port map( A1 => n4299, A2 => n4300, A3 => n4301, A4 => n4302
                           , ZN => n4298);
   U1627 : NAND4_X1 port map( A1 => n4330, A2 => n4331, A3 => n4332, A4 => 
                           n4333, ZN => n4299);
   U1628 : NAND4_X1 port map( A1 => n4321, A2 => n4322, A3 => n4323, A4 => 
                           n4324, ZN => n4300);
   U1629 : NOR2_X1 port map( A1 => n3269, A2 => n5700, ZN => N8716);
   U1630 : NOR4_X1 port map( A1 => n5701, A2 => n5702, A3 => n5703, A4 => n5704
                           , ZN => n5700);
   U1631 : NAND4_X1 port map( A1 => n5732, A2 => n5733, A3 => n5734, A4 => 
                           n5735, ZN => n5701);
   U1632 : NAND4_X1 port map( A1 => n5723, A2 => n5724, A3 => n5725, A4 => 
                           n5726, ZN => n5702);
   U1633 : NOR2_X1 port map( A1 => n3280, A2 => n4257, ZN => N8749);
   U1634 : NOR4_X1 port map( A1 => n4258, A2 => n4259, A3 => n4260, A4 => n4261
                           , ZN => n4257);
   U1635 : NAND4_X1 port map( A1 => n4289, A2 => n4290, A3 => n4291, A4 => 
                           n4292, ZN => n4258);
   U1636 : NAND4_X1 port map( A1 => n4280, A2 => n4281, A3 => n4282, A4 => 
                           n4283, ZN => n4259);
   U1637 : NOR2_X1 port map( A1 => n3269, A2 => n5659, ZN => N8717);
   U1638 : NOR4_X1 port map( A1 => n5660, A2 => n5661, A3 => n5662, A4 => n5663
                           , ZN => n5659);
   U1639 : NAND4_X1 port map( A1 => n5691, A2 => n5692, A3 => n5693, A4 => 
                           n5694, ZN => n5660);
   U1640 : NAND4_X1 port map( A1 => n5682, A2 => n5683, A3 => n5684, A4 => 
                           n5685, ZN => n5661);
   U1641 : NOR2_X1 port map( A1 => n3280, A2 => n4216, ZN => N8750);
   U1642 : NOR4_X1 port map( A1 => n4217, A2 => n4218, A3 => n4219, A4 => n4220
                           , ZN => n4216);
   U1643 : NAND4_X1 port map( A1 => n4248, A2 => n4249, A3 => n4250, A4 => 
                           n4251, ZN => n4217);
   U1644 : NAND4_X1 port map( A1 => n4239, A2 => n4240, A3 => n4241, A4 => 
                           n4242, ZN => n4218);
   U1645 : NOR2_X1 port map( A1 => n3269, A2 => n5618, ZN => N8718);
   U1646 : NOR4_X1 port map( A1 => n5619, A2 => n5620, A3 => n5621, A4 => n5622
                           , ZN => n5618);
   U1647 : NAND4_X1 port map( A1 => n5650, A2 => n5651, A3 => n5652, A4 => 
                           n5653, ZN => n5619);
   U1648 : NAND4_X1 port map( A1 => n5641, A2 => n5642, A3 => n5643, A4 => 
                           n5644, ZN => n5620);
   U1649 : NOR2_X1 port map( A1 => n3281, A2 => n4175, ZN => N8751);
   U1650 : NOR4_X1 port map( A1 => n4176, A2 => n4177, A3 => n4178, A4 => n4179
                           , ZN => n4175);
   U1651 : NAND4_X1 port map( A1 => n4207, A2 => n4208, A3 => n4209, A4 => 
                           n4210, ZN => n4176);
   U1652 : NAND4_X1 port map( A1 => n4198, A2 => n4199, A3 => n4200, A4 => 
                           n4201, ZN => n4177);
   U1653 : NOR2_X1 port map( A1 => n3270, A2 => n5577, ZN => N8719);
   U1654 : NOR4_X1 port map( A1 => n5578, A2 => n5579, A3 => n5580, A4 => n5581
                           , ZN => n5577);
   U1655 : NAND4_X1 port map( A1 => n5609, A2 => n5610, A3 => n5611, A4 => 
                           n5612, ZN => n5578);
   U1656 : NAND4_X1 port map( A1 => n5600, A2 => n5601, A3 => n5602, A4 => 
                           n5603, ZN => n5579);
   U1657 : NOR2_X1 port map( A1 => n3281, A2 => n4134, ZN => N8752);
   U1658 : NOR4_X1 port map( A1 => n4135, A2 => n4136, A3 => n4137, A4 => n4138
                           , ZN => n4134);
   U1659 : NAND4_X1 port map( A1 => n4166, A2 => n4167, A3 => n4168, A4 => 
                           n4169, ZN => n4135);
   U1660 : NAND4_X1 port map( A1 => n4157, A2 => n4158, A3 => n4159, A4 => 
                           n4160, ZN => n4136);
   U1661 : NOR2_X1 port map( A1 => n3270, A2 => n5536, ZN => N8720);
   U1662 : NOR4_X1 port map( A1 => n5537, A2 => n5538, A3 => n5539, A4 => n5540
                           , ZN => n5536);
   U1663 : NAND4_X1 port map( A1 => n5568, A2 => n5569, A3 => n5570, A4 => 
                           n5571, ZN => n5537);
   U1664 : NAND4_X1 port map( A1 => n5559, A2 => n5560, A3 => n5561, A4 => 
                           n5562, ZN => n5538);
   U1665 : NOR2_X1 port map( A1 => n3281, A2 => n4093, ZN => N8753);
   U1666 : NOR4_X1 port map( A1 => n4094, A2 => n4095, A3 => n4096, A4 => n4097
                           , ZN => n4093);
   U1667 : NAND4_X1 port map( A1 => n4125, A2 => n4126, A3 => n4127, A4 => 
                           n4128, ZN => n4094);
   U1668 : NAND4_X1 port map( A1 => n4116, A2 => n4117, A3 => n4118, A4 => 
                           n4119, ZN => n4095);
   U1669 : NOR2_X1 port map( A1 => n3270, A2 => n5495, ZN => N8721);
   U1670 : NOR4_X1 port map( A1 => n5496, A2 => n5497, A3 => n5498, A4 => n5499
                           , ZN => n5495);
   U1671 : NAND4_X1 port map( A1 => n5527, A2 => n5528, A3 => n5529, A4 => 
                           n5530, ZN => n5496);
   U1672 : NAND4_X1 port map( A1 => n5518, A2 => n5519, A3 => n5520, A4 => 
                           n5521, ZN => n5497);
   U1673 : NOR2_X1 port map( A1 => n3281, A2 => n4052, ZN => N8754);
   U1674 : NOR4_X1 port map( A1 => n4053, A2 => n4054, A3 => n4055, A4 => n4056
                           , ZN => n4052);
   U1675 : NAND4_X1 port map( A1 => n4084, A2 => n4085, A3 => n4086, A4 => 
                           n4087, ZN => n4053);
   U1676 : NAND4_X1 port map( A1 => n4075, A2 => n4076, A3 => n4077, A4 => 
                           n4078, ZN => n4054);
   U1677 : NOR2_X1 port map( A1 => n3270, A2 => n5454, ZN => N8722);
   U1678 : NOR4_X1 port map( A1 => n5455, A2 => n5456, A3 => n5457, A4 => n5458
                           , ZN => n5454);
   U1679 : NAND4_X1 port map( A1 => n5486, A2 => n5487, A3 => n5488, A4 => 
                           n5489, ZN => n5455);
   U1680 : NAND4_X1 port map( A1 => n5477, A2 => n5478, A3 => n5479, A4 => 
                           n5480, ZN => n5456);
   U1681 : NOR2_X1 port map( A1 => n3282, A2 => n4011, ZN => N8755);
   U1682 : NOR4_X1 port map( A1 => n4012, A2 => n4013, A3 => n4014, A4 => n4015
                           , ZN => n4011);
   U1683 : NAND4_X1 port map( A1 => n4043, A2 => n4044, A3 => n4045, A4 => 
                           n4046, ZN => n4012);
   U1684 : NAND4_X1 port map( A1 => n4034, A2 => n4035, A3 => n4036, A4 => 
                           n4037, ZN => n4013);
   U1685 : NOR2_X1 port map( A1 => n3272, A2 => n5413, ZN => N8723);
   U1686 : NOR4_X1 port map( A1 => n5414, A2 => n5415, A3 => n5416, A4 => n5417
                           , ZN => n5413);
   U1687 : NAND4_X1 port map( A1 => n5445, A2 => n5446, A3 => n5447, A4 => 
                           n5448, ZN => n5414);
   U1688 : NAND4_X1 port map( A1 => n5436, A2 => n5437, A3 => n5438, A4 => 
                           n5439, ZN => n5415);
   U1689 : NOR2_X1 port map( A1 => n3282, A2 => n3970, ZN => N8756);
   U1690 : NOR4_X1 port map( A1 => n3971, A2 => n3972, A3 => n3973, A4 => n3974
                           , ZN => n3970);
   U1691 : NAND4_X1 port map( A1 => n4002, A2 => n4003, A3 => n4004, A4 => 
                           n4005, ZN => n3971);
   U1692 : NAND4_X1 port map( A1 => n3993, A2 => n3994, A3 => n3995, A4 => 
                           n3996, ZN => n3972);
   U1693 : NOR2_X1 port map( A1 => n3272, A2 => n5372, ZN => N8724);
   U1694 : NOR4_X1 port map( A1 => n5373, A2 => n5374, A3 => n5375, A4 => n5376
                           , ZN => n5372);
   U1695 : NAND4_X1 port map( A1 => n5404, A2 => n5405, A3 => n5406, A4 => 
                           n5407, ZN => n5373);
   U1696 : NAND4_X1 port map( A1 => n5395, A2 => n5396, A3 => n5397, A4 => 
                           n5398, ZN => n5374);
   U1697 : NOR2_X1 port map( A1 => n3282, A2 => n3929, ZN => N8757);
   U1698 : NOR4_X1 port map( A1 => n3930, A2 => n3931, A3 => n3932, A4 => n3933
                           , ZN => n3929);
   U1699 : NAND4_X1 port map( A1 => n3961, A2 => n3962, A3 => n3963, A4 => 
                           n3964, ZN => n3930);
   U1700 : NAND4_X1 port map( A1 => n3952, A2 => n3953, A3 => n3954, A4 => 
                           n3955, ZN => n3931);
   U1701 : NOR2_X1 port map( A1 => n3272, A2 => n5331, ZN => N8725);
   U1702 : NOR4_X1 port map( A1 => n5332, A2 => n5333, A3 => n5334, A4 => n5335
                           , ZN => n5331);
   U1703 : NAND4_X1 port map( A1 => n5363, A2 => n5364, A3 => n5365, A4 => 
                           n5366, ZN => n5332);
   U1704 : NAND4_X1 port map( A1 => n5354, A2 => n5355, A3 => n5356, A4 => 
                           n5357, ZN => n5333);
   U1705 : NOR2_X1 port map( A1 => n3282, A2 => n3888, ZN => N8758);
   U1706 : NOR4_X1 port map( A1 => n3889, A2 => n3890, A3 => n3891, A4 => n3892
                           , ZN => n3888);
   U1707 : NAND4_X1 port map( A1 => n3920, A2 => n3921, A3 => n3922, A4 => 
                           n3923, ZN => n3889);
   U1708 : NAND4_X1 port map( A1 => n3911, A2 => n3912, A3 => n3913, A4 => 
                           n3914, ZN => n3890);
   U1709 : NOR2_X1 port map( A1 => n3272, A2 => n5290, ZN => N8726);
   U1710 : NOR4_X1 port map( A1 => n5291, A2 => n5292, A3 => n5293, A4 => n5294
                           , ZN => n5290);
   U1711 : NAND4_X1 port map( A1 => n5322, A2 => n5323, A3 => n5324, A4 => 
                           n5325, ZN => n5291);
   U1712 : NAND4_X1 port map( A1 => n5313, A2 => n5314, A3 => n5315, A4 => 
                           n5316, ZN => n5292);
   U1713 : NOR2_X1 port map( A1 => n3284, A2 => n3847, ZN => N8759);
   U1714 : NOR4_X1 port map( A1 => n3848, A2 => n3849, A3 => n3850, A4 => n3851
                           , ZN => n3847);
   U1715 : NAND4_X1 port map( A1 => n3879, A2 => n3880, A3 => n3881, A4 => 
                           n3882, ZN => n3848);
   U1716 : NAND4_X1 port map( A1 => n3870, A2 => n3871, A3 => n3872, A4 => 
                           n3873, ZN => n3849);
   U1717 : NOR2_X1 port map( A1 => n3273, A2 => n5249, ZN => N8727);
   U1718 : NOR4_X1 port map( A1 => n5250, A2 => n5251, A3 => n5252, A4 => n5253
                           , ZN => n5249);
   U1719 : NAND4_X1 port map( A1 => n5281, A2 => n5282, A3 => n5283, A4 => 
                           n5284, ZN => n5250);
   U1720 : NAND4_X1 port map( A1 => n5272, A2 => n5273, A3 => n5274, A4 => 
                           n5275, ZN => n5251);
   U1721 : NOR2_X1 port map( A1 => n3284, A2 => n3806, ZN => N8760);
   U1722 : NOR4_X1 port map( A1 => n3807, A2 => n3808, A3 => n3809, A4 => n3810
                           , ZN => n3806);
   U1723 : NAND4_X1 port map( A1 => n3838, A2 => n3839, A3 => n3840, A4 => 
                           n3841, ZN => n3807);
   U1724 : NAND4_X1 port map( A1 => n3829, A2 => n3830, A3 => n3831, A4 => 
                           n3832, ZN => n3808);
   U1725 : NOR2_X1 port map( A1 => n3273, A2 => n5208, ZN => N8728);
   U1726 : NOR4_X1 port map( A1 => n5209, A2 => n5210, A3 => n5211, A4 => n5212
                           , ZN => n5208);
   U1727 : NAND4_X1 port map( A1 => n5240, A2 => n5241, A3 => n5242, A4 => 
                           n5243, ZN => n5209);
   U1728 : NAND4_X1 port map( A1 => n5231, A2 => n5232, A3 => n5233, A4 => 
                           n5234, ZN => n5210);
   U1729 : NOR2_X1 port map( A1 => n3284, A2 => n3765, ZN => N8761);
   U1730 : NOR4_X1 port map( A1 => n3766, A2 => n3767, A3 => n3768, A4 => n3769
                           , ZN => n3765);
   U1731 : NAND4_X1 port map( A1 => n3797, A2 => n3798, A3 => n3799, A4 => 
                           n3800, ZN => n3766);
   U1732 : NAND4_X1 port map( A1 => n3788, A2 => n3789, A3 => n3790, A4 => 
                           n3791, ZN => n3767);
   U1733 : NOR2_X1 port map( A1 => n3273, A2 => n5167, ZN => N8729);
   U1734 : NOR4_X1 port map( A1 => n5168, A2 => n5169, A3 => n5170, A4 => n5171
                           , ZN => n5167);
   U1735 : NAND4_X1 port map( A1 => n5199, A2 => n5200, A3 => n5201, A4 => 
                           n5202, ZN => n5168);
   U1736 : NAND4_X1 port map( A1 => n5190, A2 => n5191, A3 => n5192, A4 => 
                           n5193, ZN => n5169);
   U1737 : NOR2_X1 port map( A1 => n3284, A2 => n3724, ZN => N8762);
   U1738 : NOR4_X1 port map( A1 => n3725, A2 => n3726, A3 => n3727, A4 => n3728
                           , ZN => n3724);
   U1739 : NAND4_X1 port map( A1 => n3756, A2 => n3757, A3 => n3758, A4 => 
                           n3759, ZN => n3725);
   U1740 : NAND4_X1 port map( A1 => n3747, A2 => n3748, A3 => n3749, A4 => 
                           n3750, ZN => n3726);
   U1741 : NOR2_X1 port map( A1 => n3273, A2 => n5126, ZN => N8730);
   U1742 : NOR4_X1 port map( A1 => n5127, A2 => n5128, A3 => n5129, A4 => n5130
                           , ZN => n5126);
   U1743 : NAND4_X1 port map( A1 => n5158, A2 => n5159, A3 => n5160, A4 => 
                           n5161, ZN => n5127);
   U1744 : NAND4_X1 port map( A1 => n5149, A2 => n5150, A3 => n5151, A4 => 
                           n5152, ZN => n5128);
   U1745 : NOR2_X1 port map( A1 => n3285, A2 => n3683, ZN => N8763);
   U1746 : NOR4_X1 port map( A1 => n3684, A2 => n3685, A3 => n3686, A4 => n3687
                           , ZN => n3683);
   U1747 : NAND4_X1 port map( A1 => n3715, A2 => n3716, A3 => n3717, A4 => 
                           n3718, ZN => n3684);
   U1748 : NAND4_X1 port map( A1 => n3706, A2 => n3707, A3 => n3708, A4 => 
                           n3709, ZN => n3685);
   U1749 : NOR2_X1 port map( A1 => n3274, A2 => n5085, ZN => N8731);
   U1750 : NOR4_X1 port map( A1 => n5086, A2 => n5087, A3 => n5088, A4 => n5089
                           , ZN => n5085);
   U1751 : NAND4_X1 port map( A1 => n5117, A2 => n5118, A3 => n5119, A4 => 
                           n5120, ZN => n5086);
   U1752 : NAND4_X1 port map( A1 => n5108, A2 => n5109, A3 => n5110, A4 => 
                           n5111, ZN => n5087);
   U1753 : NOR2_X1 port map( A1 => n3285, A2 => n3642, ZN => N8764);
   U1754 : NOR4_X1 port map( A1 => n3643, A2 => n3644, A3 => n3645, A4 => n3646
                           , ZN => n3642);
   U1755 : NAND4_X1 port map( A1 => n3674, A2 => n3675, A3 => n3676, A4 => 
                           n3677, ZN => n3643);
   U1756 : NAND4_X1 port map( A1 => n3665, A2 => n3666, A3 => n3667, A4 => 
                           n3668, ZN => n3644);
   U1757 : NOR2_X1 port map( A1 => n3274, A2 => n5044, ZN => N8732);
   U1758 : NOR4_X1 port map( A1 => n5045, A2 => n5046, A3 => n5047, A4 => n5048
                           , ZN => n5044);
   U1759 : NAND4_X1 port map( A1 => n5076, A2 => n5077, A3 => n5078, A4 => 
                           n5079, ZN => n5045);
   U1760 : NAND4_X1 port map( A1 => n5067, A2 => n5068, A3 => n5069, A4 => 
                           n5070, ZN => n5046);
   U1761 : NOR2_X1 port map( A1 => n3285, A2 => n3601, ZN => N8765);
   U1762 : NOR4_X1 port map( A1 => n3602, A2 => n3603, A3 => n3604, A4 => n3605
                           , ZN => n3601);
   U1763 : NAND4_X1 port map( A1 => n3633, A2 => n3634, A3 => n3635, A4 => 
                           n3636, ZN => n3602);
   U1764 : NAND4_X1 port map( A1 => n3624, A2 => n3625, A3 => n3626, A4 => 
                           n3627, ZN => n3603);
   U1765 : NOR2_X1 port map( A1 => n3274, A2 => n5003, ZN => N8733);
   U1766 : NOR4_X1 port map( A1 => n5004, A2 => n5005, A3 => n5006, A4 => n5007
                           , ZN => n5003);
   U1767 : NAND4_X1 port map( A1 => n5035, A2 => n5036, A3 => n5037, A4 => 
                           n5038, ZN => n5004);
   U1768 : NAND4_X1 port map( A1 => n5026, A2 => n5027, A3 => n5028, A4 => 
                           n5029, ZN => n5005);
   U1769 : NOR2_X1 port map( A1 => n3285, A2 => n3560, ZN => N8766);
   U1770 : NOR4_X1 port map( A1 => n3561, A2 => n3562, A3 => n3563, A4 => n3564
                           , ZN => n3560);
   U1771 : NAND4_X1 port map( A1 => n3592, A2 => n3593, A3 => n3594, A4 => 
                           n3595, ZN => n3561);
   U1772 : NAND4_X1 port map( A1 => n3583, A2 => n3584, A3 => n3585, A4 => 
                           n3586, ZN => n3562);
   U1773 : NOR2_X1 port map( A1 => n3274, A2 => n4874, ZN => N8734);
   U1774 : NOR4_X1 port map( A1 => n4875, A2 => n4876, A3 => n4877, A4 => n4878
                           , ZN => n4874);
   U1775 : NAND4_X1 port map( A1 => n4972, A2 => n4973, A3 => n4974, A4 => 
                           n4975, ZN => n4875);
   U1776 : NAND4_X1 port map( A1 => n4941, A2 => n4942, A3 => n4943, A4 => 
                           n4944, ZN => n4876);
   U1777 : NOR2_X1 port map( A1 => n3276, A2 => n3431, ZN => N8767);
   U1778 : NOR4_X1 port map( A1 => n3432, A2 => n3433, A3 => n3434, A4 => n3435
                           , ZN => n3431);
   U1779 : NAND4_X1 port map( A1 => n3529, A2 => n3530, A3 => n3531, A4 => 
                           n3532, ZN => n3432);
   U1780 : NAND4_X1 port map( A1 => n3498, A2 => n3499, A3 => n3500, A4 => 
                           n3501, ZN => n3433);
   U1781 : OAI21_X1 port map( B1 => n10920, B2 => n10921, A => n3415, ZN => 
                           n3416);
   U1782 : INV_X1 port map( A => ENABLE, ZN => n10920);
   U1783 : NAND2_X1 port map( A1 => CALL, A2 => ENABLE, ZN => n3415);
   U1784 : AND3_X1 port map( A1 => n3428, A2 => n10921, A3 => n3416, ZN => 
                           n3420);
   U1785 : NAND2_X1 port map( A1 => CWP_6_port, A2 => n3429, ZN => n3428);
   U1786 : AND3_X1 port map( A1 => n3416, A2 => n3419, A3 => RETRN, ZN => n3422
                           );
   U1787 : OAI211_X1 port map( C1 => n2898, C2 => n3416, A => n3417, B => n3418
                           , ZN => n9133);
   U1788 : OAI211_X1 port map( C1 => n3392, C2 => N8834, A => n3416, B => RETRN
                           , ZN => n3418);
   U1789 : NAND2_X1 port map( A1 => n2, A2 => n3420, ZN => n3417);
   U1790 : XNOR2_X1 port map( A => CWP_6_port, B => sub_189_carry_6_port, ZN =>
                           N8834);
   U1791 : OAI21_X1 port map( B1 => n3416, B2 => n2916, A => n3421, ZN => n9134
                           );
   U1792 : AOI22_X1 port map( A1 => N8833, A2 => n3422, B1 => n1, B2 => n3420, 
                           ZN => n3421);
   U1793 : XNOR2_X1 port map( A => CWP_5_port, B => CWP_4_port, ZN => N8833);
   U1794 : OAI21_X1 port map( B1 => n3416, B2 => N8791, A => n3423, ZN => n9135
                           );
   U1795 : AOI22_X1 port map( A1 => N8791, A2 => n3422, B1 => N8791, B2 => 
                           n3420, ZN => n3423);
   U1796 : OAI21_X1 port map( B1 => n3416, B2 => n2918, A => n3424, ZN => n9136
                           );
   U1797 : AOI22_X1 port map( A1 => N8790, A2 => n3422, B1 => N8790, B2 => 
                           n3420, ZN => n3424);
   U1798 : OAI21_X1 port map( B1 => n3416, B2 => n2919, A => n3425, ZN => n9137
                           );
   U1799 : AOI22_X1 port map( A1 => N8789, A2 => n3422, B1 => N8789, B2 => 
                           n3420, ZN => n3425);
   U1800 : OAI21_X1 port map( B1 => n3416, B2 => n2920, A => n3426, ZN => n9138
                           );
   U1801 : AOI22_X1 port map( A1 => N8788, A2 => n3422, B1 => N8788, B2 => 
                           n3420, ZN => n3426);
   U1802 : OAI21_X1 port map( B1 => n3416, B2 => n2921, A => n3427, ZN => n9139
                           );
   U1803 : AOI22_X1 port map( A1 => N8787, A2 => n3422, B1 => N8787, B2 => 
                           n3420, ZN => n3427);
   U1804 : INV_X1 port map( A => RETRN, ZN => n10921);
   U1805 : NAND2_X1 port map( A1 => n3429, A2 => n2898, ZN => n3419);
   U1806 : OR2_X1 port map( A1 => CWP_5_port, A2 => CWP_4_port, ZN => 
                           sub_189_carry_6_port);
   U1807 : AND4_X1 port map( A1 => n2920, A2 => n2919, A3 => n2921, A4 => n3430
                           , ZN => n3429);
   U1808 : NOR3_X1 port map( A1 => N8790, A2 => CWP_5_port, A3 => CWP_4_port, 
                           ZN => n3430);
   U1809 : XOR2_X1 port map( A => n2898, B => n3, Z => n2);
   U1810 : NAND2_X1 port map( A1 => CWP_5_port, A2 => CWP_4_port, ZN => n3);
   U1811 : AOI22_X1 port map( A1 => N2164, A2 => n3391, B1 => N2157, B2 => 
                           N2151, ZN => n3109);
   U1812 : XNOR2_X1 port map( A => ADD_WR(4), B => ADD_WR(3), ZN => N2164);
   U1813 : AOI22_X1 port map( A1 => N8429, A2 => n10918, B1 => N8422, B2 => 
                           N8415, ZN => n6264);
   U1814 : INV_X1 port map( A => N8430, ZN => N8429);
   U1815 : AOI22_X1 port map( A1 => N8573, A2 => n10919, B1 => N8566, B2 => 
                           N8559, ZN => n4821);
   U1816 : INV_X1 port map( A => N8574, ZN => N8573);
   U1817 : AOI22_X1 port map( A1 => ADD_RD1(2), A2 => n10918, B1 => N8419, B2 
                           => N8415, ZN => n6315);
   U1818 : AOI22_X1 port map( A1 => ADD_RD2(2), A2 => n10919, B1 => N8563, B2 
                           => N8559, ZN => n4872);
   U1819 : AOI22_X1 port map( A1 => N8428, A2 => n10918, B1 => N8421, B2 => 
                           N8415, ZN => n6265);
   U1820 : XNOR2_X1 port map( A => ADD_RD1(4), B => ADD_RD1(3), ZN => N8428);
   U1821 : AOI22_X1 port map( A1 => N8572, A2 => n10919, B1 => N8565, B2 => 
                           N8559, ZN => n4822);
   U1822 : XNOR2_X1 port map( A => ADD_RD2(4), B => ADD_RD2(3), ZN => N8572);
   U1823 : AOI22_X1 port map( A1 => ADD_RD1(1), A2 => n10918, B1 => N8418, B2 
                           => N8415, ZN => n6314);
   U1824 : AOI22_X1 port map( A1 => ADD_RD2(1), A2 => n10919, B1 => N8562, B2 
                           => N8559, ZN => n4871);
   U1825 : AOI22_X1 port map( A1 => N8427, A2 => n10918, B1 => N8420, B2 => 
                           N8415, ZN => n6280);
   U1826 : INV_X1 port map( A => ADD_RD1(3), ZN => N8427);
   U1827 : AOI22_X1 port map( A1 => N8571, A2 => n10919, B1 => N8564, B2 => 
                           N8559, ZN => n4837);
   U1828 : INV_X1 port map( A => ADD_RD2(3), ZN => N8571);
   U1829 : AOI22_X1 port map( A1 => ADD_RD1(0), A2 => n10918, B1 => N8417, B2 
                           => N8415, ZN => n6278);
   U1830 : AOI22_X1 port map( A1 => ADD_RD2(0), A2 => n10919, B1 => N8561, B2 
                           => N8559, ZN => n4835);
   U1831 : AOI222_X1 port map( A1 => n668, A2 => REGISTERS_19_0_port, B1 => 
                           n667, B2 => REGISTERS_21_0_port, C1 => n664, C2 => 
                           REGISTERS_20_0_port, ZN => n6239);
   U1832 : AOI222_X1 port map( A1 => n602, A2 => REGISTERS_41_0_port, B1 => 
                           n601, B2 => REGISTERS_43_0_port, C1 => n598, C2 => 
                           REGISTERS_42_0_port, ZN => n6270);
   U1833 : AOI222_X1 port map( A1 => n440, A2 => REGISTERS_52_0_port, B1 => 
                           n439, B2 => REGISTERS_54_0_port, C1 => n436, C2 => 
                           REGISTERS_53_0_port, ZN => n6289);
   U1834 : AOI222_X1 port map( A1 => n22, A2 => REGISTERS_85_0_port, B1 => n21,
                           B2 => REGISTERS_87_0_port, C1 => n18, C2 => 
                           REGISTERS_86_0_port, ZN => n6302);
   U1835 : AOI222_X1 port map( A1 => n1380, A2 => REGISTERS_19_0_port, B1 => 
                           n1379, B2 => REGISTERS_21_0_port, C1 => n1376, C2 =>
                           REGISTERS_20_0_port, ZN => n4796);
   U1836 : AOI222_X1 port map( A1 => n1314, A2 => REGISTERS_41_0_port, B1 => 
                           n1313, B2 => REGISTERS_43_0_port, C1 => n1310, C2 =>
                           REGISTERS_42_0_port, ZN => n4827);
   U1837 : AOI222_X1 port map( A1 => n1152, A2 => REGISTERS_52_0_port, B1 => 
                           n1151, B2 => REGISTERS_54_0_port, C1 => n1148, C2 =>
                           REGISTERS_53_0_port, ZN => n4846);
   U1838 : AOI222_X1 port map( A1 => n734, A2 => REGISTERS_85_0_port, B1 => 
                           n733, B2 => REGISTERS_87_0_port, C1 => n730, C2 => 
                           REGISTERS_86_0_port, ZN => n4859);
   U1839 : AOI222_X1 port map( A1 => n668, A2 => REGISTERS_19_1_port, B1 => 
                           n667, B2 => REGISTERS_21_1_port, C1 => n664, C2 => 
                           REGISTERS_20_1_port, ZN => n6198);
   U1840 : AOI222_X1 port map( A1 => n602, A2 => REGISTERS_41_1_port, B1 => 
                           n601, B2 => REGISTERS_43_1_port, C1 => n598, C2 => 
                           REGISTERS_42_1_port, ZN => n6207);
   U1841 : AOI222_X1 port map( A1 => n440, A2 => REGISTERS_52_1_port, B1 => 
                           n439, B2 => REGISTERS_54_1_port, C1 => n436, C2 => 
                           REGISTERS_53_1_port, ZN => n6216);
   U1842 : AOI222_X1 port map( A1 => n22, A2 => REGISTERS_85_1_port, B1 => n21,
                           B2 => REGISTERS_87_1_port, C1 => n18, C2 => 
                           REGISTERS_86_1_port, ZN => n6225);
   U1843 : AOI222_X1 port map( A1 => n1380, A2 => REGISTERS_19_1_port, B1 => 
                           n1379, B2 => REGISTERS_21_1_port, C1 => n1376, C2 =>
                           REGISTERS_20_1_port, ZN => n4755);
   U1844 : AOI222_X1 port map( A1 => n1314, A2 => REGISTERS_41_1_port, B1 => 
                           n1313, B2 => REGISTERS_43_1_port, C1 => n1310, C2 =>
                           REGISTERS_42_1_port, ZN => n4764);
   U1845 : AOI222_X1 port map( A1 => n1152, A2 => REGISTERS_52_1_port, B1 => 
                           n1151, B2 => REGISTERS_54_1_port, C1 => n1148, C2 =>
                           REGISTERS_53_1_port, ZN => n4773);
   U1846 : AOI222_X1 port map( A1 => n734, A2 => REGISTERS_85_1_port, B1 => 
                           n733, B2 => REGISTERS_87_1_port, C1 => n730, C2 => 
                           REGISTERS_86_1_port, ZN => n4782);
   U1847 : AOI222_X1 port map( A1 => n668, A2 => REGISTERS_19_2_port, B1 => 
                           n667, B2 => REGISTERS_21_2_port, C1 => n664, C2 => 
                           REGISTERS_20_2_port, ZN => n6157);
   U1848 : AOI222_X1 port map( A1 => n602, A2 => REGISTERS_41_2_port, B1 => 
                           n601, B2 => REGISTERS_43_2_port, C1 => n598, C2 => 
                           REGISTERS_42_2_port, ZN => n6166);
   U1849 : AOI222_X1 port map( A1 => n440, A2 => REGISTERS_52_2_port, B1 => 
                           n439, B2 => REGISTERS_54_2_port, C1 => n436, C2 => 
                           REGISTERS_53_2_port, ZN => n6175);
   U1850 : AOI222_X1 port map( A1 => n22, A2 => REGISTERS_85_2_port, B1 => n21,
                           B2 => REGISTERS_87_2_port, C1 => n18, C2 => 
                           REGISTERS_86_2_port, ZN => n6184);
   U1851 : AOI222_X1 port map( A1 => n1380, A2 => REGISTERS_19_2_port, B1 => 
                           n1379, B2 => REGISTERS_21_2_port, C1 => n1376, C2 =>
                           REGISTERS_20_2_port, ZN => n4714);
   U1852 : AOI222_X1 port map( A1 => n1314, A2 => REGISTERS_41_2_port, B1 => 
                           n1313, B2 => REGISTERS_43_2_port, C1 => n1310, C2 =>
                           REGISTERS_42_2_port, ZN => n4723);
   U1853 : AOI222_X1 port map( A1 => n1152, A2 => REGISTERS_52_2_port, B1 => 
                           n1151, B2 => REGISTERS_54_2_port, C1 => n1148, C2 =>
                           REGISTERS_53_2_port, ZN => n4732);
   U1854 : AOI222_X1 port map( A1 => n734, A2 => REGISTERS_85_2_port, B1 => 
                           n733, B2 => REGISTERS_87_2_port, C1 => n730, C2 => 
                           REGISTERS_86_2_port, ZN => n4741);
   U1855 : AOI222_X1 port map( A1 => n668, A2 => REGISTERS_19_3_port, B1 => 
                           n667, B2 => REGISTERS_21_3_port, C1 => n664, C2 => 
                           REGISTERS_20_3_port, ZN => n6116);
   U1856 : AOI222_X1 port map( A1 => n602, A2 => REGISTERS_41_3_port, B1 => 
                           n601, B2 => REGISTERS_43_3_port, C1 => n598, C2 => 
                           REGISTERS_42_3_port, ZN => n6125);
   U1857 : AOI222_X1 port map( A1 => n440, A2 => REGISTERS_52_3_port, B1 => 
                           n439, B2 => REGISTERS_54_3_port, C1 => n436, C2 => 
                           REGISTERS_53_3_port, ZN => n6134);
   U1858 : AOI222_X1 port map( A1 => n22, A2 => REGISTERS_85_3_port, B1 => n21,
                           B2 => REGISTERS_87_3_port, C1 => n18, C2 => 
                           REGISTERS_86_3_port, ZN => n6143);
   U1859 : AOI222_X1 port map( A1 => n1380, A2 => REGISTERS_19_3_port, B1 => 
                           n1379, B2 => REGISTERS_21_3_port, C1 => n1376, C2 =>
                           REGISTERS_20_3_port, ZN => n4673);
   U1860 : AOI222_X1 port map( A1 => n1314, A2 => REGISTERS_41_3_port, B1 => 
                           n1313, B2 => REGISTERS_43_3_port, C1 => n1310, C2 =>
                           REGISTERS_42_3_port, ZN => n4682);
   U1861 : AOI222_X1 port map( A1 => n1152, A2 => REGISTERS_52_3_port, B1 => 
                           n1151, B2 => REGISTERS_54_3_port, C1 => n1148, C2 =>
                           REGISTERS_53_3_port, ZN => n4691);
   U1862 : AOI222_X1 port map( A1 => n734, A2 => REGISTERS_85_3_port, B1 => 
                           n733, B2 => REGISTERS_87_3_port, C1 => n730, C2 => 
                           REGISTERS_86_3_port, ZN => n4700);
   U1863 : AOI222_X1 port map( A1 => n668, A2 => REGISTERS_19_4_port, B1 => 
                           n667, B2 => REGISTERS_21_4_port, C1 => n664, C2 => 
                           REGISTERS_20_4_port, ZN => n6075);
   U1864 : AOI222_X1 port map( A1 => n602, A2 => REGISTERS_41_4_port, B1 => 
                           n601, B2 => REGISTERS_43_4_port, C1 => n598, C2 => 
                           REGISTERS_42_4_port, ZN => n6084);
   U1865 : AOI222_X1 port map( A1 => n440, A2 => REGISTERS_52_4_port, B1 => 
                           n439, B2 => REGISTERS_54_4_port, C1 => n436, C2 => 
                           REGISTERS_53_4_port, ZN => n6093);
   U1866 : AOI222_X1 port map( A1 => n22, A2 => REGISTERS_85_4_port, B1 => n21,
                           B2 => REGISTERS_87_4_port, C1 => n18, C2 => 
                           REGISTERS_86_4_port, ZN => n6102);
   U1867 : AOI222_X1 port map( A1 => n1380, A2 => REGISTERS_19_4_port, B1 => 
                           n1379, B2 => REGISTERS_21_4_port, C1 => n1376, C2 =>
                           REGISTERS_20_4_port, ZN => n4632);
   U1868 : AOI222_X1 port map( A1 => n1314, A2 => REGISTERS_41_4_port, B1 => 
                           n1313, B2 => REGISTERS_43_4_port, C1 => n1310, C2 =>
                           REGISTERS_42_4_port, ZN => n4641);
   U1869 : AOI222_X1 port map( A1 => n1152, A2 => REGISTERS_52_4_port, B1 => 
                           n1151, B2 => REGISTERS_54_4_port, C1 => n1148, C2 =>
                           REGISTERS_53_4_port, ZN => n4650);
   U1870 : AOI222_X1 port map( A1 => n734, A2 => REGISTERS_85_4_port, B1 => 
                           n733, B2 => REGISTERS_87_4_port, C1 => n730, C2 => 
                           REGISTERS_86_4_port, ZN => n4659);
   U1871 : AOI222_X1 port map( A1 => n668, A2 => REGISTERS_19_5_port, B1 => 
                           n667, B2 => REGISTERS_21_5_port, C1 => n664, C2 => 
                           REGISTERS_20_5_port, ZN => n6034);
   U1872 : AOI222_X1 port map( A1 => n602, A2 => REGISTERS_41_5_port, B1 => 
                           n601, B2 => REGISTERS_43_5_port, C1 => n598, C2 => 
                           REGISTERS_42_5_port, ZN => n6043);
   U1873 : AOI222_X1 port map( A1 => n440, A2 => REGISTERS_52_5_port, B1 => 
                           n439, B2 => REGISTERS_54_5_port, C1 => n436, C2 => 
                           REGISTERS_53_5_port, ZN => n6052);
   U1874 : AOI222_X1 port map( A1 => n22, A2 => REGISTERS_85_5_port, B1 => n21,
                           B2 => REGISTERS_87_5_port, C1 => n18, C2 => 
                           REGISTERS_86_5_port, ZN => n6061);
   U1875 : AOI222_X1 port map( A1 => n1380, A2 => REGISTERS_19_5_port, B1 => 
                           n1379, B2 => REGISTERS_21_5_port, C1 => n1376, C2 =>
                           REGISTERS_20_5_port, ZN => n4591);
   U1876 : AOI222_X1 port map( A1 => n1314, A2 => REGISTERS_41_5_port, B1 => 
                           n1313, B2 => REGISTERS_43_5_port, C1 => n1310, C2 =>
                           REGISTERS_42_5_port, ZN => n4600);
   U1877 : AOI222_X1 port map( A1 => n1152, A2 => REGISTERS_52_5_port, B1 => 
                           n1151, B2 => REGISTERS_54_5_port, C1 => n1148, C2 =>
                           REGISTERS_53_5_port, ZN => n4609);
   U1878 : AOI222_X1 port map( A1 => n734, A2 => REGISTERS_85_5_port, B1 => 
                           n733, B2 => REGISTERS_87_5_port, C1 => n730, C2 => 
                           REGISTERS_86_5_port, ZN => n4618);
   U1879 : AOI222_X1 port map( A1 => n668, A2 => REGISTERS_19_6_port, B1 => 
                           n667, B2 => REGISTERS_21_6_port, C1 => n664, C2 => 
                           REGISTERS_20_6_port, ZN => n5993);
   U1880 : AOI222_X1 port map( A1 => n602, A2 => REGISTERS_41_6_port, B1 => 
                           n601, B2 => REGISTERS_43_6_port, C1 => n598, C2 => 
                           REGISTERS_42_6_port, ZN => n6002);
   U1881 : AOI222_X1 port map( A1 => n440, A2 => REGISTERS_52_6_port, B1 => 
                           n439, B2 => REGISTERS_54_6_port, C1 => n436, C2 => 
                           REGISTERS_53_6_port, ZN => n6011);
   U1882 : AOI222_X1 port map( A1 => n22, A2 => REGISTERS_85_6_port, B1 => n21,
                           B2 => REGISTERS_87_6_port, C1 => n18, C2 => 
                           REGISTERS_86_6_port, ZN => n6020);
   U1883 : AOI222_X1 port map( A1 => n1380, A2 => REGISTERS_19_6_port, B1 => 
                           n1379, B2 => REGISTERS_21_6_port, C1 => n1376, C2 =>
                           REGISTERS_20_6_port, ZN => n4550);
   U1884 : AOI222_X1 port map( A1 => n1314, A2 => REGISTERS_41_6_port, B1 => 
                           n1313, B2 => REGISTERS_43_6_port, C1 => n1310, C2 =>
                           REGISTERS_42_6_port, ZN => n4559);
   U1885 : AOI222_X1 port map( A1 => n1152, A2 => REGISTERS_52_6_port, B1 => 
                           n1151, B2 => REGISTERS_54_6_port, C1 => n1148, C2 =>
                           REGISTERS_53_6_port, ZN => n4568);
   U1886 : AOI222_X1 port map( A1 => n734, A2 => REGISTERS_85_6_port, B1 => 
                           n733, B2 => REGISTERS_87_6_port, C1 => n730, C2 => 
                           REGISTERS_86_6_port, ZN => n4577);
   U1887 : AOI222_X1 port map( A1 => n668, A2 => REGISTERS_19_7_port, B1 => 
                           n667, B2 => REGISTERS_21_7_port, C1 => n664, C2 => 
                           REGISTERS_20_7_port, ZN => n5952);
   U1888 : AOI222_X1 port map( A1 => n602, A2 => REGISTERS_41_7_port, B1 => 
                           n601, B2 => REGISTERS_43_7_port, C1 => n598, C2 => 
                           REGISTERS_42_7_port, ZN => n5961);
   U1889 : AOI222_X1 port map( A1 => n440, A2 => REGISTERS_52_7_port, B1 => 
                           n439, B2 => REGISTERS_54_7_port, C1 => n436, C2 => 
                           REGISTERS_53_7_port, ZN => n5970);
   U1890 : AOI222_X1 port map( A1 => n22, A2 => REGISTERS_85_7_port, B1 => n21,
                           B2 => REGISTERS_87_7_port, C1 => n18, C2 => 
                           REGISTERS_86_7_port, ZN => n5979);
   U1891 : AOI222_X1 port map( A1 => n1380, A2 => REGISTERS_19_7_port, B1 => 
                           n1379, B2 => REGISTERS_21_7_port, C1 => n1376, C2 =>
                           REGISTERS_20_7_port, ZN => n4509);
   U1892 : AOI222_X1 port map( A1 => n1314, A2 => REGISTERS_41_7_port, B1 => 
                           n1313, B2 => REGISTERS_43_7_port, C1 => n1310, C2 =>
                           REGISTERS_42_7_port, ZN => n4518);
   U1893 : AOI222_X1 port map( A1 => n1152, A2 => REGISTERS_52_7_port, B1 => 
                           n1151, B2 => REGISTERS_54_7_port, C1 => n1148, C2 =>
                           REGISTERS_53_7_port, ZN => n4527);
   U1894 : AOI222_X1 port map( A1 => n734, A2 => REGISTERS_85_7_port, B1 => 
                           n733, B2 => REGISTERS_87_7_port, C1 => n730, C2 => 
                           REGISTERS_86_7_port, ZN => n4536);
   U1895 : AOI222_X1 port map( A1 => n668, A2 => REGISTERS_19_8_port, B1 => 
                           n666, B2 => REGISTERS_21_8_port, C1 => n663, C2 => 
                           REGISTERS_20_8_port, ZN => n5911);
   U1896 : AOI222_X1 port map( A1 => n602, A2 => REGISTERS_41_8_port, B1 => 
                           n600, B2 => REGISTERS_43_8_port, C1 => n597, C2 => 
                           REGISTERS_42_8_port, ZN => n5920);
   U1897 : AOI222_X1 port map( A1 => n440, A2 => REGISTERS_52_8_port, B1 => 
                           n438, B2 => REGISTERS_54_8_port, C1 => n435, C2 => 
                           REGISTERS_53_8_port, ZN => n5929);
   U1898 : AOI222_X1 port map( A1 => n22, A2 => REGISTERS_85_8_port, B1 => n20,
                           B2 => REGISTERS_87_8_port, C1 => n16, C2 => 
                           REGISTERS_86_8_port, ZN => n5938);
   U1899 : AOI222_X1 port map( A1 => n1380, A2 => REGISTERS_19_8_port, B1 => 
                           n1378, B2 => REGISTERS_21_8_port, C1 => n1375, C2 =>
                           REGISTERS_20_8_port, ZN => n4468);
   U1900 : AOI222_X1 port map( A1 => n1314, A2 => REGISTERS_41_8_port, B1 => 
                           n1312, B2 => REGISTERS_43_8_port, C1 => n1309, C2 =>
                           REGISTERS_42_8_port, ZN => n4477);
   U1901 : AOI222_X1 port map( A1 => n1152, A2 => REGISTERS_52_8_port, B1 => 
                           n1150, B2 => REGISTERS_54_8_port, C1 => n1147, C2 =>
                           REGISTERS_53_8_port, ZN => n4486);
   U1902 : AOI222_X1 port map( A1 => n734, A2 => REGISTERS_85_8_port, B1 => 
                           n732, B2 => REGISTERS_87_8_port, C1 => n729, C2 => 
                           REGISTERS_86_8_port, ZN => n4495);
   U1903 : AOI222_X1 port map( A1 => n668, A2 => REGISTERS_19_9_port, B1 => 
                           n666, B2 => REGISTERS_21_9_port, C1 => n663, C2 => 
                           REGISTERS_20_9_port, ZN => n5870);
   U1904 : AOI222_X1 port map( A1 => n602, A2 => REGISTERS_41_9_port, B1 => 
                           n600, B2 => REGISTERS_43_9_port, C1 => n597, C2 => 
                           REGISTERS_42_9_port, ZN => n5879);
   U1905 : AOI222_X1 port map( A1 => n440, A2 => REGISTERS_52_9_port, B1 => 
                           n438, B2 => REGISTERS_54_9_port, C1 => n435, C2 => 
                           REGISTERS_53_9_port, ZN => n5888);
   U1906 : AOI222_X1 port map( A1 => n22, A2 => REGISTERS_85_9_port, B1 => n20,
                           B2 => REGISTERS_87_9_port, C1 => n16, C2 => 
                           REGISTERS_86_9_port, ZN => n5897);
   U1907 : AOI222_X1 port map( A1 => n1380, A2 => REGISTERS_19_9_port, B1 => 
                           n1378, B2 => REGISTERS_21_9_port, C1 => n1375, C2 =>
                           REGISTERS_20_9_port, ZN => n4427);
   U1908 : AOI222_X1 port map( A1 => n1314, A2 => REGISTERS_41_9_port, B1 => 
                           n1312, B2 => REGISTERS_43_9_port, C1 => n1309, C2 =>
                           REGISTERS_42_9_port, ZN => n4436);
   U1909 : AOI222_X1 port map( A1 => n1152, A2 => REGISTERS_52_9_port, B1 => 
                           n1150, B2 => REGISTERS_54_9_port, C1 => n1147, C2 =>
                           REGISTERS_53_9_port, ZN => n4445);
   U1910 : AOI222_X1 port map( A1 => n734, A2 => REGISTERS_85_9_port, B1 => 
                           n732, B2 => REGISTERS_87_9_port, C1 => n729, C2 => 
                           REGISTERS_86_9_port, ZN => n4454);
   U1911 : AOI222_X1 port map( A1 => n668, A2 => REGISTERS_19_10_port, B1 => 
                           n666, B2 => REGISTERS_21_10_port, C1 => n663, C2 => 
                           REGISTERS_20_10_port, ZN => n5829);
   U1912 : AOI222_X1 port map( A1 => n602, A2 => REGISTERS_41_10_port, B1 => 
                           n600, B2 => REGISTERS_43_10_port, C1 => n597, C2 => 
                           REGISTERS_42_10_port, ZN => n5838);
   U1913 : AOI222_X1 port map( A1 => n440, A2 => REGISTERS_52_10_port, B1 => 
                           n438, B2 => REGISTERS_54_10_port, C1 => n435, C2 => 
                           REGISTERS_53_10_port, ZN => n5847);
   U1914 : AOI222_X1 port map( A1 => n22, A2 => REGISTERS_85_10_port, B1 => n20
                           , B2 => REGISTERS_87_10_port, C1 => n16, C2 => 
                           REGISTERS_86_10_port, ZN => n5856);
   U1915 : AOI222_X1 port map( A1 => n1380, A2 => REGISTERS_19_10_port, B1 => 
                           n1378, B2 => REGISTERS_21_10_port, C1 => n1375, C2 
                           => REGISTERS_20_10_port, ZN => n4386);
   U1916 : AOI222_X1 port map( A1 => n1314, A2 => REGISTERS_41_10_port, B1 => 
                           n1312, B2 => REGISTERS_43_10_port, C1 => n1309, C2 
                           => REGISTERS_42_10_port, ZN => n4395);
   U1917 : AOI222_X1 port map( A1 => n1152, A2 => REGISTERS_52_10_port, B1 => 
                           n1150, B2 => REGISTERS_54_10_port, C1 => n1147, C2 
                           => REGISTERS_53_10_port, ZN => n4404);
   U1918 : AOI222_X1 port map( A1 => n734, A2 => REGISTERS_85_10_port, B1 => 
                           n732, B2 => REGISTERS_87_10_port, C1 => n729, C2 => 
                           REGISTERS_86_10_port, ZN => n4413);
   U1919 : AOI222_X1 port map( A1 => n668, A2 => REGISTERS_19_11_port, B1 => 
                           n666, B2 => REGISTERS_21_11_port, C1 => n663, C2 => 
                           REGISTERS_20_11_port, ZN => n5788);
   U1920 : AOI222_X1 port map( A1 => n602, A2 => REGISTERS_41_11_port, B1 => 
                           n600, B2 => REGISTERS_43_11_port, C1 => n597, C2 => 
                           REGISTERS_42_11_port, ZN => n5797);
   U1921 : AOI222_X1 port map( A1 => n440, A2 => REGISTERS_52_11_port, B1 => 
                           n438, B2 => REGISTERS_54_11_port, C1 => n435, C2 => 
                           REGISTERS_53_11_port, ZN => n5806);
   U1922 : AOI222_X1 port map( A1 => n22, A2 => REGISTERS_85_11_port, B1 => n20
                           , B2 => REGISTERS_87_11_port, C1 => n16, C2 => 
                           REGISTERS_86_11_port, ZN => n5815);
   U1923 : AOI222_X1 port map( A1 => n1380, A2 => REGISTERS_19_11_port, B1 => 
                           n1378, B2 => REGISTERS_21_11_port, C1 => n1375, C2 
                           => REGISTERS_20_11_port, ZN => n4345);
   U1924 : AOI222_X1 port map( A1 => n1314, A2 => REGISTERS_41_11_port, B1 => 
                           n1312, B2 => REGISTERS_43_11_port, C1 => n1309, C2 
                           => REGISTERS_42_11_port, ZN => n4354);
   U1925 : AOI222_X1 port map( A1 => n1152, A2 => REGISTERS_52_11_port, B1 => 
                           n1150, B2 => REGISTERS_54_11_port, C1 => n1147, C2 
                           => REGISTERS_53_11_port, ZN => n4363);
   U1926 : AOI222_X1 port map( A1 => n734, A2 => REGISTERS_85_11_port, B1 => 
                           n732, B2 => REGISTERS_87_11_port, C1 => n729, C2 => 
                           REGISTERS_86_11_port, ZN => n4372);
   U1927 : AOI222_X1 port map( A1 => n669, A2 => REGISTERS_19_12_port, B1 => 
                           n666, B2 => REGISTERS_21_12_port, C1 => n663, C2 => 
                           REGISTERS_20_12_port, ZN => n5747);
   U1928 : AOI222_X1 port map( A1 => n603, A2 => REGISTERS_41_12_port, B1 => 
                           n600, B2 => REGISTERS_43_12_port, C1 => n597, C2 => 
                           REGISTERS_42_12_port, ZN => n5756);
   U1929 : AOI222_X1 port map( A1 => n441, A2 => REGISTERS_52_12_port, B1 => 
                           n438, B2 => REGISTERS_54_12_port, C1 => n435, C2 => 
                           REGISTERS_53_12_port, ZN => n5765);
   U1930 : AOI222_X1 port map( A1 => n23, A2 => REGISTERS_85_12_port, B1 => n20
                           , B2 => REGISTERS_87_12_port, C1 => n16, C2 => 
                           REGISTERS_86_12_port, ZN => n5774);
   U1931 : AOI222_X1 port map( A1 => n1381, A2 => REGISTERS_19_12_port, B1 => 
                           n1378, B2 => REGISTERS_21_12_port, C1 => n1375, C2 
                           => REGISTERS_20_12_port, ZN => n4304);
   U1932 : AOI222_X1 port map( A1 => n1315, A2 => REGISTERS_41_12_port, B1 => 
                           n1312, B2 => REGISTERS_43_12_port, C1 => n1309, C2 
                           => REGISTERS_42_12_port, ZN => n4313);
   U1933 : AOI222_X1 port map( A1 => n1153, A2 => REGISTERS_52_12_port, B1 => 
                           n1150, B2 => REGISTERS_54_12_port, C1 => n1147, C2 
                           => REGISTERS_53_12_port, ZN => n4322);
   U1934 : AOI222_X1 port map( A1 => n735, A2 => REGISTERS_85_12_port, B1 => 
                           n732, B2 => REGISTERS_87_12_port, C1 => n729, C2 => 
                           REGISTERS_86_12_port, ZN => n4331);
   U1935 : AOI222_X1 port map( A1 => n669, A2 => REGISTERS_19_13_port, B1 => 
                           n666, B2 => REGISTERS_21_13_port, C1 => n663, C2 => 
                           REGISTERS_20_13_port, ZN => n5706);
   U1936 : AOI222_X1 port map( A1 => n603, A2 => REGISTERS_41_13_port, B1 => 
                           n600, B2 => REGISTERS_43_13_port, C1 => n597, C2 => 
                           REGISTERS_42_13_port, ZN => n5715);
   U1937 : AOI222_X1 port map( A1 => n441, A2 => REGISTERS_52_13_port, B1 => 
                           n438, B2 => REGISTERS_54_13_port, C1 => n435, C2 => 
                           REGISTERS_53_13_port, ZN => n5724);
   U1938 : AOI222_X1 port map( A1 => n23, A2 => REGISTERS_85_13_port, B1 => n20
                           , B2 => REGISTERS_87_13_port, C1 => n16, C2 => 
                           REGISTERS_86_13_port, ZN => n5733);
   U1939 : AOI222_X1 port map( A1 => n1381, A2 => REGISTERS_19_13_port, B1 => 
                           n1378, B2 => REGISTERS_21_13_port, C1 => n1375, C2 
                           => REGISTERS_20_13_port, ZN => n4263);
   U1940 : AOI222_X1 port map( A1 => n1315, A2 => REGISTERS_41_13_port, B1 => 
                           n1312, B2 => REGISTERS_43_13_port, C1 => n1309, C2 
                           => REGISTERS_42_13_port, ZN => n4272);
   U1941 : AOI222_X1 port map( A1 => n1153, A2 => REGISTERS_52_13_port, B1 => 
                           n1150, B2 => REGISTERS_54_13_port, C1 => n1147, C2 
                           => REGISTERS_53_13_port, ZN => n4281);
   U1942 : AOI222_X1 port map( A1 => n735, A2 => REGISTERS_85_13_port, B1 => 
                           n732, B2 => REGISTERS_87_13_port, C1 => n729, C2 => 
                           REGISTERS_86_13_port, ZN => n4290);
   U1943 : AOI222_X1 port map( A1 => n669, A2 => REGISTERS_19_14_port, B1 => 
                           n666, B2 => REGISTERS_21_14_port, C1 => n663, C2 => 
                           REGISTERS_20_14_port, ZN => n5665);
   U1944 : AOI222_X1 port map( A1 => n603, A2 => REGISTERS_41_14_port, B1 => 
                           n600, B2 => REGISTERS_43_14_port, C1 => n597, C2 => 
                           REGISTERS_42_14_port, ZN => n5674);
   U1945 : AOI222_X1 port map( A1 => n441, A2 => REGISTERS_52_14_port, B1 => 
                           n438, B2 => REGISTERS_54_14_port, C1 => n435, C2 => 
                           REGISTERS_53_14_port, ZN => n5683);
   U1946 : AOI222_X1 port map( A1 => n23, A2 => REGISTERS_85_14_port, B1 => n20
                           , B2 => REGISTERS_87_14_port, C1 => n16, C2 => 
                           REGISTERS_86_14_port, ZN => n5692);
   U1947 : AOI222_X1 port map( A1 => n1381, A2 => REGISTERS_19_14_port, B1 => 
                           n1378, B2 => REGISTERS_21_14_port, C1 => n1375, C2 
                           => REGISTERS_20_14_port, ZN => n4222);
   U1948 : AOI222_X1 port map( A1 => n1315, A2 => REGISTERS_41_14_port, B1 => 
                           n1312, B2 => REGISTERS_43_14_port, C1 => n1309, C2 
                           => REGISTERS_42_14_port, ZN => n4231);
   U1949 : AOI222_X1 port map( A1 => n1153, A2 => REGISTERS_52_14_port, B1 => 
                           n1150, B2 => REGISTERS_54_14_port, C1 => n1147, C2 
                           => REGISTERS_53_14_port, ZN => n4240);
   U1950 : AOI222_X1 port map( A1 => n735, A2 => REGISTERS_85_14_port, B1 => 
                           n732, B2 => REGISTERS_87_14_port, C1 => n729, C2 => 
                           REGISTERS_86_14_port, ZN => n4249);
   U1951 : AOI222_X1 port map( A1 => n669, A2 => REGISTERS_19_15_port, B1 => 
                           n666, B2 => REGISTERS_21_15_port, C1 => n663, C2 => 
                           REGISTERS_20_15_port, ZN => n5624);
   U1952 : AOI222_X1 port map( A1 => n603, A2 => REGISTERS_41_15_port, B1 => 
                           n600, B2 => REGISTERS_43_15_port, C1 => n597, C2 => 
                           REGISTERS_42_15_port, ZN => n5633);
   U1953 : AOI222_X1 port map( A1 => n441, A2 => REGISTERS_52_15_port, B1 => 
                           n438, B2 => REGISTERS_54_15_port, C1 => n435, C2 => 
                           REGISTERS_53_15_port, ZN => n5642);
   U1954 : AOI222_X1 port map( A1 => n23, A2 => REGISTERS_85_15_port, B1 => n20
                           , B2 => REGISTERS_87_15_port, C1 => n16, C2 => 
                           REGISTERS_86_15_port, ZN => n5651);
   U1955 : AOI222_X1 port map( A1 => n1381, A2 => REGISTERS_19_15_port, B1 => 
                           n1378, B2 => REGISTERS_21_15_port, C1 => n1375, C2 
                           => REGISTERS_20_15_port, ZN => n4181);
   U1956 : AOI222_X1 port map( A1 => n1315, A2 => REGISTERS_41_15_port, B1 => 
                           n1312, B2 => REGISTERS_43_15_port, C1 => n1309, C2 
                           => REGISTERS_42_15_port, ZN => n4190);
   U1957 : AOI222_X1 port map( A1 => n1153, A2 => REGISTERS_52_15_port, B1 => 
                           n1150, B2 => REGISTERS_54_15_port, C1 => n1147, C2 
                           => REGISTERS_53_15_port, ZN => n4199);
   U1958 : AOI222_X1 port map( A1 => n735, A2 => REGISTERS_85_15_port, B1 => 
                           n732, B2 => REGISTERS_87_15_port, C1 => n729, C2 => 
                           REGISTERS_86_15_port, ZN => n4208);
   U1959 : AOI222_X1 port map( A1 => n669, A2 => REGISTERS_19_16_port, B1 => 
                           n666, B2 => REGISTERS_21_16_port, C1 => n663, C2 => 
                           REGISTERS_20_16_port, ZN => n5583);
   U1960 : AOI222_X1 port map( A1 => n603, A2 => REGISTERS_41_16_port, B1 => 
                           n600, B2 => REGISTERS_43_16_port, C1 => n597, C2 => 
                           REGISTERS_42_16_port, ZN => n5592);
   U1961 : AOI222_X1 port map( A1 => n441, A2 => REGISTERS_52_16_port, B1 => 
                           n438, B2 => REGISTERS_54_16_port, C1 => n435, C2 => 
                           REGISTERS_53_16_port, ZN => n5601);
   U1962 : AOI222_X1 port map( A1 => n23, A2 => REGISTERS_85_16_port, B1 => n20
                           , B2 => REGISTERS_87_16_port, C1 => n16, C2 => 
                           REGISTERS_86_16_port, ZN => n5610);
   U1963 : AOI222_X1 port map( A1 => n1381, A2 => REGISTERS_19_16_port, B1 => 
                           n1378, B2 => REGISTERS_21_16_port, C1 => n1375, C2 
                           => REGISTERS_20_16_port, ZN => n4140);
   U1964 : AOI222_X1 port map( A1 => n1315, A2 => REGISTERS_41_16_port, B1 => 
                           n1312, B2 => REGISTERS_43_16_port, C1 => n1309, C2 
                           => REGISTERS_42_16_port, ZN => n4149);
   U1965 : AOI222_X1 port map( A1 => n1153, A2 => REGISTERS_52_16_port, B1 => 
                           n1150, B2 => REGISTERS_54_16_port, C1 => n1147, C2 
                           => REGISTERS_53_16_port, ZN => n4158);
   U1966 : AOI222_X1 port map( A1 => n735, A2 => REGISTERS_85_16_port, B1 => 
                           n732, B2 => REGISTERS_87_16_port, C1 => n729, C2 => 
                           REGISTERS_86_16_port, ZN => n4167);
   U1967 : AOI222_X1 port map( A1 => n669, A2 => REGISTERS_19_17_port, B1 => 
                           n666, B2 => REGISTERS_21_17_port, C1 => n663, C2 => 
                           REGISTERS_20_17_port, ZN => n5542);
   U1968 : AOI222_X1 port map( A1 => n603, A2 => REGISTERS_41_17_port, B1 => 
                           n600, B2 => REGISTERS_43_17_port, C1 => n597, C2 => 
                           REGISTERS_42_17_port, ZN => n5551);
   U1969 : AOI222_X1 port map( A1 => n441, A2 => REGISTERS_52_17_port, B1 => 
                           n438, B2 => REGISTERS_54_17_port, C1 => n435, C2 => 
                           REGISTERS_53_17_port, ZN => n5560);
   U1970 : AOI222_X1 port map( A1 => n23, A2 => REGISTERS_85_17_port, B1 => n20
                           , B2 => REGISTERS_87_17_port, C1 => n16, C2 => 
                           REGISTERS_86_17_port, ZN => n5569);
   U1971 : AOI222_X1 port map( A1 => n1381, A2 => REGISTERS_19_17_port, B1 => 
                           n1378, B2 => REGISTERS_21_17_port, C1 => n1375, C2 
                           => REGISTERS_20_17_port, ZN => n4099);
   U1972 : AOI222_X1 port map( A1 => n1315, A2 => REGISTERS_41_17_port, B1 => 
                           n1312, B2 => REGISTERS_43_17_port, C1 => n1309, C2 
                           => REGISTERS_42_17_port, ZN => n4108);
   U1973 : AOI222_X1 port map( A1 => n1153, A2 => REGISTERS_52_17_port, B1 => 
                           n1150, B2 => REGISTERS_54_17_port, C1 => n1147, C2 
                           => REGISTERS_53_17_port, ZN => n4117);
   U1974 : AOI222_X1 port map( A1 => n735, A2 => REGISTERS_85_17_port, B1 => 
                           n732, B2 => REGISTERS_87_17_port, C1 => n729, C2 => 
                           REGISTERS_86_17_port, ZN => n4126);
   U1975 : AOI222_X1 port map( A1 => n669, A2 => REGISTERS_19_18_port, B1 => 
                           n666, B2 => REGISTERS_21_18_port, C1 => n663, C2 => 
                           REGISTERS_20_18_port, ZN => n5501);
   U1976 : AOI222_X1 port map( A1 => n603, A2 => REGISTERS_41_18_port, B1 => 
                           n600, B2 => REGISTERS_43_18_port, C1 => n597, C2 => 
                           REGISTERS_42_18_port, ZN => n5510);
   U1977 : AOI222_X1 port map( A1 => n441, A2 => REGISTERS_52_18_port, B1 => 
                           n438, B2 => REGISTERS_54_18_port, C1 => n435, C2 => 
                           REGISTERS_53_18_port, ZN => n5519);
   U1978 : AOI222_X1 port map( A1 => n23, A2 => REGISTERS_85_18_port, B1 => n20
                           , B2 => REGISTERS_87_18_port, C1 => n16, C2 => 
                           REGISTERS_86_18_port, ZN => n5528);
   U1979 : AOI222_X1 port map( A1 => n1381, A2 => REGISTERS_19_18_port, B1 => 
                           n1378, B2 => REGISTERS_21_18_port, C1 => n1375, C2 
                           => REGISTERS_20_18_port, ZN => n4058);
   U1980 : AOI222_X1 port map( A1 => n1315, A2 => REGISTERS_41_18_port, B1 => 
                           n1312, B2 => REGISTERS_43_18_port, C1 => n1309, C2 
                           => REGISTERS_42_18_port, ZN => n4067);
   U1981 : AOI222_X1 port map( A1 => n1153, A2 => REGISTERS_52_18_port, B1 => 
                           n1150, B2 => REGISTERS_54_18_port, C1 => n1147, C2 
                           => REGISTERS_53_18_port, ZN => n4076);
   U1982 : AOI222_X1 port map( A1 => n735, A2 => REGISTERS_85_18_port, B1 => 
                           n732, B2 => REGISTERS_87_18_port, C1 => n729, C2 => 
                           REGISTERS_86_18_port, ZN => n4085);
   U1983 : AOI222_X1 port map( A1 => n669, A2 => REGISTERS_19_19_port, B1 => 
                           n666, B2 => REGISTERS_21_19_port, C1 => n663, C2 => 
                           REGISTERS_20_19_port, ZN => n5460);
   U1984 : AOI222_X1 port map( A1 => n603, A2 => REGISTERS_41_19_port, B1 => 
                           n600, B2 => REGISTERS_43_19_port, C1 => n597, C2 => 
                           REGISTERS_42_19_port, ZN => n5469);
   U1985 : AOI222_X1 port map( A1 => n441, A2 => REGISTERS_52_19_port, B1 => 
                           n438, B2 => REGISTERS_54_19_port, C1 => n435, C2 => 
                           REGISTERS_53_19_port, ZN => n5478);
   U1986 : AOI222_X1 port map( A1 => n23, A2 => REGISTERS_85_19_port, B1 => n20
                           , B2 => REGISTERS_87_19_port, C1 => n16, C2 => 
                           REGISTERS_86_19_port, ZN => n5487);
   U1987 : AOI222_X1 port map( A1 => n1381, A2 => REGISTERS_19_19_port, B1 => 
                           n1378, B2 => REGISTERS_21_19_port, C1 => n1375, C2 
                           => REGISTERS_20_19_port, ZN => n4017);
   U1988 : AOI222_X1 port map( A1 => n1315, A2 => REGISTERS_41_19_port, B1 => 
                           n1312, B2 => REGISTERS_43_19_port, C1 => n1309, C2 
                           => REGISTERS_42_19_port, ZN => n4026);
   U1989 : AOI222_X1 port map( A1 => n1153, A2 => REGISTERS_52_19_port, B1 => 
                           n1150, B2 => REGISTERS_54_19_port, C1 => n1147, C2 
                           => REGISTERS_53_19_port, ZN => n4035);
   U1990 : AOI222_X1 port map( A1 => n735, A2 => REGISTERS_85_19_port, B1 => 
                           n732, B2 => REGISTERS_87_19_port, C1 => n729, C2 => 
                           REGISTERS_86_19_port, ZN => n4044);
   U1991 : AOI222_X1 port map( A1 => n669, A2 => REGISTERS_19_20_port, B1 => 
                           n665, B2 => REGISTERS_21_20_port, C1 => n662, C2 => 
                           REGISTERS_20_20_port, ZN => n5419);
   U1992 : AOI222_X1 port map( A1 => n603, A2 => REGISTERS_41_20_port, B1 => 
                           n599, B2 => REGISTERS_43_20_port, C1 => n596, C2 => 
                           REGISTERS_42_20_port, ZN => n5428);
   U1993 : AOI222_X1 port map( A1 => n441, A2 => REGISTERS_52_20_port, B1 => 
                           n437, B2 => REGISTERS_54_20_port, C1 => n434, C2 => 
                           REGISTERS_53_20_port, ZN => n5437);
   U1994 : AOI222_X1 port map( A1 => n23, A2 => REGISTERS_85_20_port, B1 => n19
                           , B2 => REGISTERS_87_20_port, C1 => n15, C2 => 
                           REGISTERS_86_20_port, ZN => n5446);
   U1995 : AOI222_X1 port map( A1 => n1381, A2 => REGISTERS_19_20_port, B1 => 
                           n1377, B2 => REGISTERS_21_20_port, C1 => n1374, C2 
                           => REGISTERS_20_20_port, ZN => n3976);
   U1996 : AOI222_X1 port map( A1 => n1315, A2 => REGISTERS_41_20_port, B1 => 
                           n1311, B2 => REGISTERS_43_20_port, C1 => n1308, C2 
                           => REGISTERS_42_20_port, ZN => n3985);
   U1997 : AOI222_X1 port map( A1 => n1153, A2 => REGISTERS_52_20_port, B1 => 
                           n1149, B2 => REGISTERS_54_20_port, C1 => n1146, C2 
                           => REGISTERS_53_20_port, ZN => n3994);
   U1998 : AOI222_X1 port map( A1 => n735, A2 => REGISTERS_85_20_port, B1 => 
                           n731, B2 => REGISTERS_87_20_port, C1 => n728, C2 => 
                           REGISTERS_86_20_port, ZN => n4003);
   U1999 : AOI222_X1 port map( A1 => n669, A2 => REGISTERS_19_21_port, B1 => 
                           n665, B2 => REGISTERS_21_21_port, C1 => n662, C2 => 
                           REGISTERS_20_21_port, ZN => n5378);
   U2000 : AOI222_X1 port map( A1 => n603, A2 => REGISTERS_41_21_port, B1 => 
                           n599, B2 => REGISTERS_43_21_port, C1 => n596, C2 => 
                           REGISTERS_42_21_port, ZN => n5387);
   U2001 : AOI222_X1 port map( A1 => n441, A2 => REGISTERS_52_21_port, B1 => 
                           n437, B2 => REGISTERS_54_21_port, C1 => n434, C2 => 
                           REGISTERS_53_21_port, ZN => n5396);
   U2002 : AOI222_X1 port map( A1 => n23, A2 => REGISTERS_85_21_port, B1 => n19
                           , B2 => REGISTERS_87_21_port, C1 => n15, C2 => 
                           REGISTERS_86_21_port, ZN => n5405);
   U2003 : AOI222_X1 port map( A1 => n1381, A2 => REGISTERS_19_21_port, B1 => 
                           n1377, B2 => REGISTERS_21_21_port, C1 => n1374, C2 
                           => REGISTERS_20_21_port, ZN => n3935);
   U2004 : AOI222_X1 port map( A1 => n1315, A2 => REGISTERS_41_21_port, B1 => 
                           n1311, B2 => REGISTERS_43_21_port, C1 => n1308, C2 
                           => REGISTERS_42_21_port, ZN => n3944);
   U2005 : AOI222_X1 port map( A1 => n1153, A2 => REGISTERS_52_21_port, B1 => 
                           n1149, B2 => REGISTERS_54_21_port, C1 => n1146, C2 
                           => REGISTERS_53_21_port, ZN => n3953);
   U2006 : AOI222_X1 port map( A1 => n735, A2 => REGISTERS_85_21_port, B1 => 
                           n731, B2 => REGISTERS_87_21_port, C1 => n728, C2 => 
                           REGISTERS_86_21_port, ZN => n3962);
   U2007 : AOI222_X1 port map( A1 => n669, A2 => REGISTERS_19_22_port, B1 => 
                           n665, B2 => REGISTERS_21_22_port, C1 => n662, C2 => 
                           REGISTERS_20_22_port, ZN => n5337);
   U2008 : AOI222_X1 port map( A1 => n603, A2 => REGISTERS_41_22_port, B1 => 
                           n599, B2 => REGISTERS_43_22_port, C1 => n596, C2 => 
                           REGISTERS_42_22_port, ZN => n5346);
   U2009 : AOI222_X1 port map( A1 => n441, A2 => REGISTERS_52_22_port, B1 => 
                           n437, B2 => REGISTERS_54_22_port, C1 => n434, C2 => 
                           REGISTERS_53_22_port, ZN => n5355);
   U2010 : AOI222_X1 port map( A1 => n23, A2 => REGISTERS_85_22_port, B1 => n19
                           , B2 => REGISTERS_87_22_port, C1 => n15, C2 => 
                           REGISTERS_86_22_port, ZN => n5364);
   U2011 : AOI222_X1 port map( A1 => n1381, A2 => REGISTERS_19_22_port, B1 => 
                           n1377, B2 => REGISTERS_21_22_port, C1 => n1374, C2 
                           => REGISTERS_20_22_port, ZN => n3894);
   U2012 : AOI222_X1 port map( A1 => n1315, A2 => REGISTERS_41_22_port, B1 => 
                           n1311, B2 => REGISTERS_43_22_port, C1 => n1308, C2 
                           => REGISTERS_42_22_port, ZN => n3903);
   U2013 : AOI222_X1 port map( A1 => n1153, A2 => REGISTERS_52_22_port, B1 => 
                           n1149, B2 => REGISTERS_54_22_port, C1 => n1146, C2 
                           => REGISTERS_53_22_port, ZN => n3912);
   U2014 : AOI222_X1 port map( A1 => n735, A2 => REGISTERS_85_22_port, B1 => 
                           n731, B2 => REGISTERS_87_22_port, C1 => n728, C2 => 
                           REGISTERS_86_22_port, ZN => n3921);
   U2015 : AOI222_X1 port map( A1 => n669, A2 => REGISTERS_19_23_port, B1 => 
                           n665, B2 => REGISTERS_21_23_port, C1 => n662, C2 => 
                           REGISTERS_20_23_port, ZN => n5296);
   U2016 : AOI222_X1 port map( A1 => n603, A2 => REGISTERS_41_23_port, B1 => 
                           n599, B2 => REGISTERS_43_23_port, C1 => n596, C2 => 
                           REGISTERS_42_23_port, ZN => n5305);
   U2017 : AOI222_X1 port map( A1 => n441, A2 => REGISTERS_52_23_port, B1 => 
                           n437, B2 => REGISTERS_54_23_port, C1 => n434, C2 => 
                           REGISTERS_53_23_port, ZN => n5314);
   U2018 : AOI222_X1 port map( A1 => n23, A2 => REGISTERS_85_23_port, B1 => n19
                           , B2 => REGISTERS_87_23_port, C1 => n15, C2 => 
                           REGISTERS_86_23_port, ZN => n5323);
   U2019 : AOI222_X1 port map( A1 => n1381, A2 => REGISTERS_19_23_port, B1 => 
                           n1377, B2 => REGISTERS_21_23_port, C1 => n1374, C2 
                           => REGISTERS_20_23_port, ZN => n3853);
   U2020 : AOI222_X1 port map( A1 => n1315, A2 => REGISTERS_41_23_port, B1 => 
                           n1311, B2 => REGISTERS_43_23_port, C1 => n1308, C2 
                           => REGISTERS_42_23_port, ZN => n3862);
   U2021 : AOI222_X1 port map( A1 => n1153, A2 => REGISTERS_52_23_port, B1 => 
                           n1149, B2 => REGISTERS_54_23_port, C1 => n1146, C2 
                           => REGISTERS_53_23_port, ZN => n3871);
   U2022 : AOI222_X1 port map( A1 => n735, A2 => REGISTERS_85_23_port, B1 => 
                           n731, B2 => REGISTERS_87_23_port, C1 => n728, C2 => 
                           REGISTERS_86_23_port, ZN => n3880);
   U2023 : AOI222_X1 port map( A1 => n670, A2 => REGISTERS_19_24_port, B1 => 
                           n665, B2 => REGISTERS_21_24_port, C1 => n662, C2 => 
                           REGISTERS_20_24_port, ZN => n5255);
   U2024 : AOI222_X1 port map( A1 => n604, A2 => REGISTERS_41_24_port, B1 => 
                           n599, B2 => REGISTERS_43_24_port, C1 => n596, C2 => 
                           REGISTERS_42_24_port, ZN => n5264);
   U2025 : AOI222_X1 port map( A1 => n442, A2 => REGISTERS_52_24_port, B1 => 
                           n437, B2 => REGISTERS_54_24_port, C1 => n434, C2 => 
                           REGISTERS_53_24_port, ZN => n5273);
   U2026 : AOI222_X1 port map( A1 => n24, A2 => REGISTERS_85_24_port, B1 => n19
                           , B2 => REGISTERS_87_24_port, C1 => n15, C2 => 
                           REGISTERS_86_24_port, ZN => n5282);
   U2027 : AOI222_X1 port map( A1 => n1382, A2 => REGISTERS_19_24_port, B1 => 
                           n1377, B2 => REGISTERS_21_24_port, C1 => n1374, C2 
                           => REGISTERS_20_24_port, ZN => n3812);
   U2028 : AOI222_X1 port map( A1 => n1316, A2 => REGISTERS_41_24_port, B1 => 
                           n1311, B2 => REGISTERS_43_24_port, C1 => n1308, C2 
                           => REGISTERS_42_24_port, ZN => n3821);
   U2029 : AOI222_X1 port map( A1 => n1154, A2 => REGISTERS_52_24_port, B1 => 
                           n1149, B2 => REGISTERS_54_24_port, C1 => n1146, C2 
                           => REGISTERS_53_24_port, ZN => n3830);
   U2030 : AOI222_X1 port map( A1 => n736, A2 => REGISTERS_85_24_port, B1 => 
                           n731, B2 => REGISTERS_87_24_port, C1 => n728, C2 => 
                           REGISTERS_86_24_port, ZN => n3839);
   U2031 : AOI222_X1 port map( A1 => n670, A2 => REGISTERS_19_25_port, B1 => 
                           n665, B2 => REGISTERS_21_25_port, C1 => n662, C2 => 
                           REGISTERS_20_25_port, ZN => n5214);
   U2032 : AOI222_X1 port map( A1 => n604, A2 => REGISTERS_41_25_port, B1 => 
                           n599, B2 => REGISTERS_43_25_port, C1 => n596, C2 => 
                           REGISTERS_42_25_port, ZN => n5223);
   U2033 : AOI222_X1 port map( A1 => n442, A2 => REGISTERS_52_25_port, B1 => 
                           n437, B2 => REGISTERS_54_25_port, C1 => n434, C2 => 
                           REGISTERS_53_25_port, ZN => n5232);
   U2034 : AOI222_X1 port map( A1 => n24, A2 => REGISTERS_85_25_port, B1 => n19
                           , B2 => REGISTERS_87_25_port, C1 => n15, C2 => 
                           REGISTERS_86_25_port, ZN => n5241);
   U2035 : AOI222_X1 port map( A1 => n1382, A2 => REGISTERS_19_25_port, B1 => 
                           n1377, B2 => REGISTERS_21_25_port, C1 => n1374, C2 
                           => REGISTERS_20_25_port, ZN => n3771);
   U2036 : AOI222_X1 port map( A1 => n1316, A2 => REGISTERS_41_25_port, B1 => 
                           n1311, B2 => REGISTERS_43_25_port, C1 => n1308, C2 
                           => REGISTERS_42_25_port, ZN => n3780);
   U2037 : AOI222_X1 port map( A1 => n1154, A2 => REGISTERS_52_25_port, B1 => 
                           n1149, B2 => REGISTERS_54_25_port, C1 => n1146, C2 
                           => REGISTERS_53_25_port, ZN => n3789);
   U2038 : AOI222_X1 port map( A1 => n736, A2 => REGISTERS_85_25_port, B1 => 
                           n731, B2 => REGISTERS_87_25_port, C1 => n728, C2 => 
                           REGISTERS_86_25_port, ZN => n3798);
   U2039 : AOI222_X1 port map( A1 => n670, A2 => REGISTERS_19_26_port, B1 => 
                           n665, B2 => REGISTERS_21_26_port, C1 => n662, C2 => 
                           REGISTERS_20_26_port, ZN => n5173);
   U2040 : AOI222_X1 port map( A1 => n604, A2 => REGISTERS_41_26_port, B1 => 
                           n599, B2 => REGISTERS_43_26_port, C1 => n596, C2 => 
                           REGISTERS_42_26_port, ZN => n5182);
   U2041 : AOI222_X1 port map( A1 => n442, A2 => REGISTERS_52_26_port, B1 => 
                           n437, B2 => REGISTERS_54_26_port, C1 => n434, C2 => 
                           REGISTERS_53_26_port, ZN => n5191);
   U2042 : AOI222_X1 port map( A1 => n24, A2 => REGISTERS_85_26_port, B1 => n19
                           , B2 => REGISTERS_87_26_port, C1 => n15, C2 => 
                           REGISTERS_86_26_port, ZN => n5200);
   U2043 : AOI222_X1 port map( A1 => n1382, A2 => REGISTERS_19_26_port, B1 => 
                           n1377, B2 => REGISTERS_21_26_port, C1 => n1374, C2 
                           => REGISTERS_20_26_port, ZN => n3730);
   U2044 : AOI222_X1 port map( A1 => n1316, A2 => REGISTERS_41_26_port, B1 => 
                           n1311, B2 => REGISTERS_43_26_port, C1 => n1308, C2 
                           => REGISTERS_42_26_port, ZN => n3739);
   U2045 : AOI222_X1 port map( A1 => n1154, A2 => REGISTERS_52_26_port, B1 => 
                           n1149, B2 => REGISTERS_54_26_port, C1 => n1146, C2 
                           => REGISTERS_53_26_port, ZN => n3748);
   U2046 : AOI222_X1 port map( A1 => n736, A2 => REGISTERS_85_26_port, B1 => 
                           n731, B2 => REGISTERS_87_26_port, C1 => n728, C2 => 
                           REGISTERS_86_26_port, ZN => n3757);
   U2047 : AOI222_X1 port map( A1 => n670, A2 => REGISTERS_19_27_port, B1 => 
                           n665, B2 => REGISTERS_21_27_port, C1 => n662, C2 => 
                           REGISTERS_20_27_port, ZN => n5132);
   U2048 : AOI222_X1 port map( A1 => n604, A2 => REGISTERS_41_27_port, B1 => 
                           n599, B2 => REGISTERS_43_27_port, C1 => n596, C2 => 
                           REGISTERS_42_27_port, ZN => n5141);
   U2049 : AOI222_X1 port map( A1 => n442, A2 => REGISTERS_52_27_port, B1 => 
                           n437, B2 => REGISTERS_54_27_port, C1 => n434, C2 => 
                           REGISTERS_53_27_port, ZN => n5150);
   U2050 : AOI222_X1 port map( A1 => n24, A2 => REGISTERS_85_27_port, B1 => n19
                           , B2 => REGISTERS_87_27_port, C1 => n15, C2 => 
                           REGISTERS_86_27_port, ZN => n5159);
   U2051 : AOI222_X1 port map( A1 => n1382, A2 => REGISTERS_19_27_port, B1 => 
                           n1377, B2 => REGISTERS_21_27_port, C1 => n1374, C2 
                           => REGISTERS_20_27_port, ZN => n3689);
   U2052 : AOI222_X1 port map( A1 => n1316, A2 => REGISTERS_41_27_port, B1 => 
                           n1311, B2 => REGISTERS_43_27_port, C1 => n1308, C2 
                           => REGISTERS_42_27_port, ZN => n3698);
   U2053 : AOI222_X1 port map( A1 => n1154, A2 => REGISTERS_52_27_port, B1 => 
                           n1149, B2 => REGISTERS_54_27_port, C1 => n1146, C2 
                           => REGISTERS_53_27_port, ZN => n3707);
   U2054 : AOI222_X1 port map( A1 => n736, A2 => REGISTERS_85_27_port, B1 => 
                           n731, B2 => REGISTERS_87_27_port, C1 => n728, C2 => 
                           REGISTERS_86_27_port, ZN => n3716);
   U2055 : AOI222_X1 port map( A1 => n670, A2 => REGISTERS_19_28_port, B1 => 
                           n665, B2 => REGISTERS_21_28_port, C1 => n662, C2 => 
                           REGISTERS_20_28_port, ZN => n5091);
   U2056 : AOI222_X1 port map( A1 => n604, A2 => REGISTERS_41_28_port, B1 => 
                           n599, B2 => REGISTERS_43_28_port, C1 => n596, C2 => 
                           REGISTERS_42_28_port, ZN => n5100);
   U2057 : AOI222_X1 port map( A1 => n442, A2 => REGISTERS_52_28_port, B1 => 
                           n437, B2 => REGISTERS_54_28_port, C1 => n434, C2 => 
                           REGISTERS_53_28_port, ZN => n5109);
   U2058 : AOI222_X1 port map( A1 => n24, A2 => REGISTERS_85_28_port, B1 => n19
                           , B2 => REGISTERS_87_28_port, C1 => n15, C2 => 
                           REGISTERS_86_28_port, ZN => n5118);
   U2059 : AOI222_X1 port map( A1 => n1382, A2 => REGISTERS_19_28_port, B1 => 
                           n1377, B2 => REGISTERS_21_28_port, C1 => n1374, C2 
                           => REGISTERS_20_28_port, ZN => n3648);
   U2060 : AOI222_X1 port map( A1 => n1316, A2 => REGISTERS_41_28_port, B1 => 
                           n1311, B2 => REGISTERS_43_28_port, C1 => n1308, C2 
                           => REGISTERS_42_28_port, ZN => n3657);
   U2061 : AOI222_X1 port map( A1 => n1154, A2 => REGISTERS_52_28_port, B1 => 
                           n1149, B2 => REGISTERS_54_28_port, C1 => n1146, C2 
                           => REGISTERS_53_28_port, ZN => n3666);
   U2062 : AOI222_X1 port map( A1 => n736, A2 => REGISTERS_85_28_port, B1 => 
                           n731, B2 => REGISTERS_87_28_port, C1 => n728, C2 => 
                           REGISTERS_86_28_port, ZN => n3675);
   U2063 : AOI222_X1 port map( A1 => n670, A2 => REGISTERS_19_29_port, B1 => 
                           n665, B2 => REGISTERS_21_29_port, C1 => n662, C2 => 
                           REGISTERS_20_29_port, ZN => n5050);
   U2064 : AOI222_X1 port map( A1 => n604, A2 => REGISTERS_41_29_port, B1 => 
                           n599, B2 => REGISTERS_43_29_port, C1 => n596, C2 => 
                           REGISTERS_42_29_port, ZN => n5059);
   U2065 : AOI222_X1 port map( A1 => n442, A2 => REGISTERS_52_29_port, B1 => 
                           n437, B2 => REGISTERS_54_29_port, C1 => n434, C2 => 
                           REGISTERS_53_29_port, ZN => n5068);
   U2066 : AOI222_X1 port map( A1 => n24, A2 => REGISTERS_85_29_port, B1 => n19
                           , B2 => REGISTERS_87_29_port, C1 => n15, C2 => 
                           REGISTERS_86_29_port, ZN => n5077);
   U2067 : AOI222_X1 port map( A1 => n1382, A2 => REGISTERS_19_29_port, B1 => 
                           n1377, B2 => REGISTERS_21_29_port, C1 => n1374, C2 
                           => REGISTERS_20_29_port, ZN => n3607);
   U2068 : AOI222_X1 port map( A1 => n1316, A2 => REGISTERS_41_29_port, B1 => 
                           n1311, B2 => REGISTERS_43_29_port, C1 => n1308, C2 
                           => REGISTERS_42_29_port, ZN => n3616);
   U2069 : AOI222_X1 port map( A1 => n1154, A2 => REGISTERS_52_29_port, B1 => 
                           n1149, B2 => REGISTERS_54_29_port, C1 => n1146, C2 
                           => REGISTERS_53_29_port, ZN => n3625);
   U2070 : AOI222_X1 port map( A1 => n736, A2 => REGISTERS_85_29_port, B1 => 
                           n731, B2 => REGISTERS_87_29_port, C1 => n728, C2 => 
                           REGISTERS_86_29_port, ZN => n3634);
   U2071 : AOI222_X1 port map( A1 => n670, A2 => REGISTERS_19_30_port, B1 => 
                           n665, B2 => REGISTERS_21_30_port, C1 => n662, C2 => 
                           REGISTERS_20_30_port, ZN => n5009);
   U2072 : AOI222_X1 port map( A1 => n604, A2 => REGISTERS_41_30_port, B1 => 
                           n599, B2 => REGISTERS_43_30_port, C1 => n596, C2 => 
                           REGISTERS_42_30_port, ZN => n5018);
   U2073 : AOI222_X1 port map( A1 => n442, A2 => REGISTERS_52_30_port, B1 => 
                           n437, B2 => REGISTERS_54_30_port, C1 => n434, C2 => 
                           REGISTERS_53_30_port, ZN => n5027);
   U2074 : AOI222_X1 port map( A1 => n24, A2 => REGISTERS_85_30_port, B1 => n19
                           , B2 => REGISTERS_87_30_port, C1 => n15, C2 => 
                           REGISTERS_86_30_port, ZN => n5036);
   U2075 : AOI222_X1 port map( A1 => n1382, A2 => REGISTERS_19_30_port, B1 => 
                           n1377, B2 => REGISTERS_21_30_port, C1 => n1374, C2 
                           => REGISTERS_20_30_port, ZN => n3566);
   U2076 : AOI222_X1 port map( A1 => n1316, A2 => REGISTERS_41_30_port, B1 => 
                           n1311, B2 => REGISTERS_43_30_port, C1 => n1308, C2 
                           => REGISTERS_42_30_port, ZN => n3575);
   U2077 : AOI222_X1 port map( A1 => n1154, A2 => REGISTERS_52_30_port, B1 => 
                           n1149, B2 => REGISTERS_54_30_port, C1 => n1146, C2 
                           => REGISTERS_53_30_port, ZN => n3584);
   U2078 : AOI222_X1 port map( A1 => n736, A2 => REGISTERS_85_30_port, B1 => 
                           n731, B2 => REGISTERS_87_30_port, C1 => n728, C2 => 
                           REGISTERS_86_30_port, ZN => n3593);
   U2079 : AOI222_X1 port map( A1 => n670, A2 => REGISTERS_19_31_port, B1 => 
                           n665, B2 => REGISTERS_21_31_port, C1 => n662, C2 => 
                           REGISTERS_20_31_port, ZN => n4880);
   U2080 : AOI222_X1 port map( A1 => n604, A2 => REGISTERS_41_31_port, B1 => 
                           n599, B2 => REGISTERS_43_31_port, C1 => n596, C2 => 
                           REGISTERS_42_31_port, ZN => n4911);
   U2081 : AOI222_X1 port map( A1 => n442, A2 => REGISTERS_52_31_port, B1 => 
                           n437, B2 => REGISTERS_54_31_port, C1 => n434, C2 => 
                           REGISTERS_53_31_port, ZN => n4942);
   U2082 : AOI222_X1 port map( A1 => n24, A2 => REGISTERS_85_31_port, B1 => n19
                           , B2 => REGISTERS_87_31_port, C1 => n15, C2 => 
                           REGISTERS_86_31_port, ZN => n4973);
   U2083 : AOI222_X1 port map( A1 => n1382, A2 => REGISTERS_19_31_port, B1 => 
                           n1377, B2 => REGISTERS_21_31_port, C1 => n1374, C2 
                           => REGISTERS_20_31_port, ZN => n3437);
   U2084 : AOI222_X1 port map( A1 => n1316, A2 => REGISTERS_41_31_port, B1 => 
                           n1311, B2 => REGISTERS_43_31_port, C1 => n1308, C2 
                           => REGISTERS_42_31_port, ZN => n3468);
   U2085 : AOI222_X1 port map( A1 => n1154, A2 => REGISTERS_52_31_port, B1 => 
                           n1149, B2 => REGISTERS_54_31_port, C1 => n1146, C2 
                           => REGISTERS_53_31_port, ZN => n3499);
   U2086 : AOI222_X1 port map( A1 => n736, A2 => REGISTERS_85_31_port, B1 => 
                           n731, B2 => REGISTERS_87_31_port, C1 => n728, C2 => 
                           REGISTERS_86_31_port, ZN => n3530);
   U2087 : OAI222_X1 port map( A1 => n207, A2 => n710, B1 => n239, B2 => n707, 
                           C1 => n175, C2 => n704, ZN => n6244);
   U2088 : OAI222_X1 port map( A1 => n911, A2 => n644, B1 => n943, B2 => n641, 
                           C1 => n879, C2 => n638, ZN => n6275);
   U2089 : OAI222_X1 port map( A1 => n1967, A2 => n482, B1 => n1999, B2 => n479
                           , C1 => n1935, C2 => n476, ZN => n6294);
   U2090 : OAI222_X1 port map( A1 => n2319, A2 => n64, B1 => n2351, B2 => n61, 
                           C1 => n2287, C2 => n58, ZN => n6307);
   U2091 : OAI222_X1 port map( A1 => n207, A2 => n1422, B1 => n239, B2 => n1419
                           , C1 => n175, C2 => n1416, ZN => n4801);
   U2092 : OAI222_X1 port map( A1 => n911, A2 => n1356, B1 => n943, B2 => n1353
                           , C1 => n879, C2 => n1350, ZN => n4832);
   U2093 : OAI222_X1 port map( A1 => n1967, A2 => n1194, B1 => n1999, B2 => 
                           n1191, C1 => n1935, C2 => n1188, ZN => n4851);
   U2094 : OAI222_X1 port map( A1 => n2319, A2 => n776, B1 => n2351, B2 => n773
                           , C1 => n2287, C2 => n770, ZN => n4864);
   U2095 : OAI222_X1 port map( A1 => n206, A2 => n710, B1 => n238, B2 => n707, 
                           C1 => n174, C2 => n704, ZN => n6203);
   U2096 : OAI222_X1 port map( A1 => n910, A2 => n644, B1 => n942, B2 => n641, 
                           C1 => n878, C2 => n638, ZN => n6212);
   U2097 : OAI222_X1 port map( A1 => n1966, A2 => n482, B1 => n1998, B2 => n479
                           , C1 => n1934, C2 => n476, ZN => n6221);
   U2098 : OAI222_X1 port map( A1 => n2318, A2 => n64, B1 => n2350, B2 => n61, 
                           C1 => n2286, C2 => n58, ZN => n6230);
   U2099 : OAI222_X1 port map( A1 => n206, A2 => n1422, B1 => n238, B2 => n1419
                           , C1 => n174, C2 => n1416, ZN => n4760);
   U2100 : OAI222_X1 port map( A1 => n910, A2 => n1356, B1 => n942, B2 => n1353
                           , C1 => n878, C2 => n1350, ZN => n4769);
   U2101 : OAI222_X1 port map( A1 => n1966, A2 => n1194, B1 => n1998, B2 => 
                           n1191, C1 => n1934, C2 => n1188, ZN => n4778);
   U2102 : OAI222_X1 port map( A1 => n2318, A2 => n776, B1 => n2350, B2 => n773
                           , C1 => n2286, C2 => n770, ZN => n4787);
   U2103 : OAI222_X1 port map( A1 => n205, A2 => n710, B1 => n237, B2 => n707, 
                           C1 => n173, C2 => n704, ZN => n6162);
   U2104 : OAI222_X1 port map( A1 => n909, A2 => n644, B1 => n941, B2 => n641, 
                           C1 => n877, C2 => n638, ZN => n6171);
   U2105 : OAI222_X1 port map( A1 => n1965, A2 => n482, B1 => n1997, B2 => n479
                           , C1 => n1933, C2 => n476, ZN => n6180);
   U2106 : OAI222_X1 port map( A1 => n2317, A2 => n64, B1 => n2349, B2 => n61, 
                           C1 => n2285, C2 => n58, ZN => n6189);
   U2107 : OAI222_X1 port map( A1 => n205, A2 => n1422, B1 => n237, B2 => n1419
                           , C1 => n173, C2 => n1416, ZN => n4719);
   U2108 : OAI222_X1 port map( A1 => n909, A2 => n1356, B1 => n941, B2 => n1353
                           , C1 => n877, C2 => n1350, ZN => n4728);
   U2109 : OAI222_X1 port map( A1 => n1965, A2 => n1194, B1 => n1997, B2 => 
                           n1191, C1 => n1933, C2 => n1188, ZN => n4737);
   U2110 : OAI222_X1 port map( A1 => n2317, A2 => n776, B1 => n2349, B2 => n773
                           , C1 => n2285, C2 => n770, ZN => n4746);
   U2111 : OAI222_X1 port map( A1 => n204, A2 => n710, B1 => n236, B2 => n707, 
                           C1 => n172, C2 => n704, ZN => n6121);
   U2112 : OAI222_X1 port map( A1 => n908, A2 => n644, B1 => n940, B2 => n641, 
                           C1 => n876, C2 => n638, ZN => n6130);
   U2113 : OAI222_X1 port map( A1 => n1964, A2 => n482, B1 => n1996, B2 => n479
                           , C1 => n1932, C2 => n476, ZN => n6139);
   U2114 : OAI222_X1 port map( A1 => n2316, A2 => n64, B1 => n2348, B2 => n61, 
                           C1 => n2284, C2 => n58, ZN => n6148);
   U2115 : OAI222_X1 port map( A1 => n204, A2 => n1422, B1 => n236, B2 => n1419
                           , C1 => n172, C2 => n1416, ZN => n4678);
   U2116 : OAI222_X1 port map( A1 => n908, A2 => n1356, B1 => n940, B2 => n1353
                           , C1 => n876, C2 => n1350, ZN => n4687);
   U2117 : OAI222_X1 port map( A1 => n1964, A2 => n1194, B1 => n1996, B2 => 
                           n1191, C1 => n1932, C2 => n1188, ZN => n4696);
   U2118 : OAI222_X1 port map( A1 => n2316, A2 => n776, B1 => n2348, B2 => n773
                           , C1 => n2284, C2 => n770, ZN => n4705);
   U2119 : OAI222_X1 port map( A1 => n203, A2 => n710, B1 => n235, B2 => n707, 
                           C1 => n171, C2 => n704, ZN => n6080);
   U2120 : OAI222_X1 port map( A1 => n907, A2 => n644, B1 => n939, B2 => n641, 
                           C1 => n875, C2 => n638, ZN => n6089);
   U2121 : OAI222_X1 port map( A1 => n1963, A2 => n482, B1 => n1995, B2 => n479
                           , C1 => n1931, C2 => n476, ZN => n6098);
   U2122 : OAI222_X1 port map( A1 => n2315, A2 => n64, B1 => n2347, B2 => n61, 
                           C1 => n2283, C2 => n58, ZN => n6107);
   U2123 : OAI222_X1 port map( A1 => n203, A2 => n1422, B1 => n235, B2 => n1419
                           , C1 => n171, C2 => n1416, ZN => n4637);
   U2124 : OAI222_X1 port map( A1 => n907, A2 => n1356, B1 => n939, B2 => n1353
                           , C1 => n875, C2 => n1350, ZN => n4646);
   U2125 : OAI222_X1 port map( A1 => n1963, A2 => n1194, B1 => n1995, B2 => 
                           n1191, C1 => n1931, C2 => n1188, ZN => n4655);
   U2126 : OAI222_X1 port map( A1 => n2315, A2 => n776, B1 => n2347, B2 => n773
                           , C1 => n2283, C2 => n770, ZN => n4664);
   U2127 : OAI222_X1 port map( A1 => n202, A2 => n710, B1 => n234, B2 => n707, 
                           C1 => n170, C2 => n704, ZN => n6039);
   U2128 : OAI222_X1 port map( A1 => n906, A2 => n644, B1 => n938, B2 => n641, 
                           C1 => n874, C2 => n638, ZN => n6048);
   U2129 : OAI222_X1 port map( A1 => n1962, A2 => n482, B1 => n1994, B2 => n479
                           , C1 => n1930, C2 => n476, ZN => n6057);
   U2130 : OAI222_X1 port map( A1 => n2314, A2 => n64, B1 => n2346, B2 => n61, 
                           C1 => n2282, C2 => n58, ZN => n6066);
   U2131 : OAI222_X1 port map( A1 => n202, A2 => n1422, B1 => n234, B2 => n1419
                           , C1 => n170, C2 => n1416, ZN => n4596);
   U2132 : OAI222_X1 port map( A1 => n906, A2 => n1356, B1 => n938, B2 => n1353
                           , C1 => n874, C2 => n1350, ZN => n4605);
   U2133 : OAI222_X1 port map( A1 => n1962, A2 => n1194, B1 => n1994, B2 => 
                           n1191, C1 => n1930, C2 => n1188, ZN => n4614);
   U2134 : OAI222_X1 port map( A1 => n2314, A2 => n776, B1 => n2346, B2 => n773
                           , C1 => n2282, C2 => n770, ZN => n4623);
   U2135 : OAI222_X1 port map( A1 => n201, A2 => n710, B1 => n233, B2 => n707, 
                           C1 => n169, C2 => n704, ZN => n5998);
   U2136 : OAI222_X1 port map( A1 => n905, A2 => n644, B1 => n937, B2 => n641, 
                           C1 => n873, C2 => n638, ZN => n6007);
   U2137 : OAI222_X1 port map( A1 => n1961, A2 => n482, B1 => n1993, B2 => n479
                           , C1 => n1929, C2 => n476, ZN => n6016);
   U2138 : OAI222_X1 port map( A1 => n2313, A2 => n64, B1 => n2345, B2 => n61, 
                           C1 => n2281, C2 => n58, ZN => n6025);
   U2139 : OAI222_X1 port map( A1 => n201, A2 => n1422, B1 => n233, B2 => n1419
                           , C1 => n169, C2 => n1416, ZN => n4555);
   U2140 : OAI222_X1 port map( A1 => n905, A2 => n1356, B1 => n937, B2 => n1353
                           , C1 => n873, C2 => n1350, ZN => n4564);
   U2141 : OAI222_X1 port map( A1 => n1961, A2 => n1194, B1 => n1993, B2 => 
                           n1191, C1 => n1929, C2 => n1188, ZN => n4573);
   U2142 : OAI222_X1 port map( A1 => n2313, A2 => n776, B1 => n2345, B2 => n773
                           , C1 => n2281, C2 => n770, ZN => n4582);
   U2143 : OAI222_X1 port map( A1 => n200, A2 => n710, B1 => n232, B2 => n707, 
                           C1 => n168, C2 => n704, ZN => n5957);
   U2144 : OAI222_X1 port map( A1 => n904, A2 => n644, B1 => n936, B2 => n641, 
                           C1 => n872, C2 => n638, ZN => n5966);
   U2145 : OAI222_X1 port map( A1 => n1960, A2 => n482, B1 => n1992, B2 => n479
                           , C1 => n1928, C2 => n476, ZN => n5975);
   U2146 : OAI222_X1 port map( A1 => n2312, A2 => n64, B1 => n2344, B2 => n61, 
                           C1 => n2280, C2 => n58, ZN => n5984);
   U2147 : OAI222_X1 port map( A1 => n200, A2 => n1422, B1 => n232, B2 => n1419
                           , C1 => n168, C2 => n1416, ZN => n4514);
   U2148 : OAI222_X1 port map( A1 => n904, A2 => n1356, B1 => n936, B2 => n1353
                           , C1 => n872, C2 => n1350, ZN => n4523);
   U2149 : OAI222_X1 port map( A1 => n1960, A2 => n1194, B1 => n1992, B2 => 
                           n1191, C1 => n1928, C2 => n1188, ZN => n4532);
   U2150 : OAI222_X1 port map( A1 => n2312, A2 => n776, B1 => n2344, B2 => n773
                           , C1 => n2280, C2 => n770, ZN => n4541);
   U2151 : OAI222_X1 port map( A1 => n199, A2 => n710, B1 => n231, B2 => n707, 
                           C1 => n167, C2 => n704, ZN => n5916);
   U2152 : OAI222_X1 port map( A1 => n903, A2 => n644, B1 => n935, B2 => n641, 
                           C1 => n871, C2 => n638, ZN => n5925);
   U2153 : OAI222_X1 port map( A1 => n1959, A2 => n482, B1 => n1991, B2 => n479
                           , C1 => n1927, C2 => n476, ZN => n5934);
   U2154 : OAI222_X1 port map( A1 => n2311, A2 => n64, B1 => n2343, B2 => n61, 
                           C1 => n2279, C2 => n58, ZN => n5943);
   U2155 : OAI222_X1 port map( A1 => n199, A2 => n1422, B1 => n231, B2 => n1419
                           , C1 => n167, C2 => n1416, ZN => n4473);
   U2156 : OAI222_X1 port map( A1 => n903, A2 => n1356, B1 => n935, B2 => n1353
                           , C1 => n871, C2 => n1350, ZN => n4482);
   U2157 : OAI222_X1 port map( A1 => n1959, A2 => n1194, B1 => n1991, B2 => 
                           n1191, C1 => n1927, C2 => n1188, ZN => n4491);
   U2158 : OAI222_X1 port map( A1 => n2311, A2 => n776, B1 => n2343, B2 => n773
                           , C1 => n2279, C2 => n770, ZN => n4500);
   U2159 : OAI222_X1 port map( A1 => n198, A2 => n710, B1 => n230, B2 => n707, 
                           C1 => n166, C2 => n704, ZN => n5875);
   U2160 : OAI222_X1 port map( A1 => n902, A2 => n644, B1 => n934, B2 => n641, 
                           C1 => n870, C2 => n638, ZN => n5884);
   U2161 : OAI222_X1 port map( A1 => n1958, A2 => n482, B1 => n1990, B2 => n479
                           , C1 => n1926, C2 => n476, ZN => n5893);
   U2162 : OAI222_X1 port map( A1 => n2310, A2 => n64, B1 => n2342, B2 => n61, 
                           C1 => n2278, C2 => n58, ZN => n5902);
   U2163 : OAI222_X1 port map( A1 => n198, A2 => n1422, B1 => n230, B2 => n1419
                           , C1 => n166, C2 => n1416, ZN => n4432);
   U2164 : OAI222_X1 port map( A1 => n902, A2 => n1356, B1 => n934, B2 => n1353
                           , C1 => n870, C2 => n1350, ZN => n4441);
   U2165 : OAI222_X1 port map( A1 => n1958, A2 => n1194, B1 => n1990, B2 => 
                           n1191, C1 => n1926, C2 => n1188, ZN => n4450);
   U2166 : OAI222_X1 port map( A1 => n2310, A2 => n776, B1 => n2342, B2 => n773
                           , C1 => n2278, C2 => n770, ZN => n4459);
   U2167 : OAI222_X1 port map( A1 => n197, A2 => n710, B1 => n229, B2 => n707, 
                           C1 => n165, C2 => n704, ZN => n5834);
   U2168 : OAI222_X1 port map( A1 => n901, A2 => n644, B1 => n933, B2 => n641, 
                           C1 => n869, C2 => n638, ZN => n5843);
   U2169 : OAI222_X1 port map( A1 => n1957, A2 => n482, B1 => n1989, B2 => n479
                           , C1 => n1925, C2 => n476, ZN => n5852);
   U2170 : OAI222_X1 port map( A1 => n2309, A2 => n64, B1 => n2341, B2 => n61, 
                           C1 => n2277, C2 => n58, ZN => n5861);
   U2171 : OAI222_X1 port map( A1 => n197, A2 => n1422, B1 => n229, B2 => n1419
                           , C1 => n165, C2 => n1416, ZN => n4391);
   U2172 : OAI222_X1 port map( A1 => n901, A2 => n1356, B1 => n933, B2 => n1353
                           , C1 => n869, C2 => n1350, ZN => n4400);
   U2173 : OAI222_X1 port map( A1 => n1957, A2 => n1194, B1 => n1989, B2 => 
                           n1191, C1 => n1925, C2 => n1188, ZN => n4409);
   U2174 : OAI222_X1 port map( A1 => n2309, A2 => n776, B1 => n2341, B2 => n773
                           , C1 => n2277, C2 => n770, ZN => n4418);
   U2175 : OAI222_X1 port map( A1 => n196, A2 => n710, B1 => n228, B2 => n707, 
                           C1 => n164, C2 => n704, ZN => n5793);
   U2176 : OAI222_X1 port map( A1 => n900, A2 => n644, B1 => n932, B2 => n641, 
                           C1 => n868, C2 => n638, ZN => n5802);
   U2177 : OAI222_X1 port map( A1 => n1956, A2 => n482, B1 => n1988, B2 => n479
                           , C1 => n1924, C2 => n476, ZN => n5811);
   U2178 : OAI222_X1 port map( A1 => n2308, A2 => n64, B1 => n2340, B2 => n61, 
                           C1 => n2276, C2 => n58, ZN => n5820);
   U2179 : OAI222_X1 port map( A1 => n196, A2 => n1422, B1 => n228, B2 => n1419
                           , C1 => n164, C2 => n1416, ZN => n4350);
   U2180 : OAI222_X1 port map( A1 => n900, A2 => n1356, B1 => n932, B2 => n1353
                           , C1 => n868, C2 => n1350, ZN => n4359);
   U2181 : OAI222_X1 port map( A1 => n1956, A2 => n1194, B1 => n1988, B2 => 
                           n1191, C1 => n1924, C2 => n1188, ZN => n4368);
   U2182 : OAI222_X1 port map( A1 => n2308, A2 => n776, B1 => n2340, B2 => n773
                           , C1 => n2276, C2 => n770, ZN => n4377);
   U2183 : OAI222_X1 port map( A1 => n195, A2 => n711, B1 => n227, B2 => n708, 
                           C1 => n163, C2 => n705, ZN => n5752);
   U2184 : OAI222_X1 port map( A1 => n899, A2 => n645, B1 => n931, B2 => n642, 
                           C1 => n867, C2 => n639, ZN => n5761);
   U2185 : OAI222_X1 port map( A1 => n1955, A2 => n483, B1 => n1987, B2 => n480
                           , C1 => n1923, C2 => n477, ZN => n5770);
   U2186 : OAI222_X1 port map( A1 => n2307, A2 => n65, B1 => n2339, B2 => n62, 
                           C1 => n2275, C2 => n59, ZN => n5779);
   U2187 : OAI222_X1 port map( A1 => n195, A2 => n1423, B1 => n227, B2 => n1420
                           , C1 => n163, C2 => n1417, ZN => n4309);
   U2188 : OAI222_X1 port map( A1 => n899, A2 => n1357, B1 => n931, B2 => n1354
                           , C1 => n867, C2 => n1351, ZN => n4318);
   U2189 : OAI222_X1 port map( A1 => n1955, A2 => n1195, B1 => n1987, B2 => 
                           n1192, C1 => n1923, C2 => n1189, ZN => n4327);
   U2190 : OAI222_X1 port map( A1 => n2307, A2 => n777, B1 => n2339, B2 => n774
                           , C1 => n2275, C2 => n771, ZN => n4336);
   U2191 : OAI222_X1 port map( A1 => n194, A2 => n711, B1 => n226, B2 => n708, 
                           C1 => n162, C2 => n705, ZN => n5711);
   U2192 : OAI222_X1 port map( A1 => n898, A2 => n645, B1 => n930, B2 => n642, 
                           C1 => n866, C2 => n639, ZN => n5720);
   U2193 : OAI222_X1 port map( A1 => n1954, A2 => n483, B1 => n1986, B2 => n480
                           , C1 => n1922, C2 => n477, ZN => n5729);
   U2194 : OAI222_X1 port map( A1 => n2306, A2 => n65, B1 => n2338, B2 => n62, 
                           C1 => n2274, C2 => n59, ZN => n5738);
   U2195 : OAI222_X1 port map( A1 => n194, A2 => n1423, B1 => n226, B2 => n1420
                           , C1 => n162, C2 => n1417, ZN => n4268);
   U2196 : OAI222_X1 port map( A1 => n898, A2 => n1357, B1 => n930, B2 => n1354
                           , C1 => n866, C2 => n1351, ZN => n4277);
   U2197 : OAI222_X1 port map( A1 => n1954, A2 => n1195, B1 => n1986, B2 => 
                           n1192, C1 => n1922, C2 => n1189, ZN => n4286);
   U2198 : OAI222_X1 port map( A1 => n2306, A2 => n777, B1 => n2338, B2 => n774
                           , C1 => n2274, C2 => n771, ZN => n4295);
   U2199 : OAI222_X1 port map( A1 => n193, A2 => n711, B1 => n225, B2 => n708, 
                           C1 => n161, C2 => n705, ZN => n5670);
   U2200 : OAI222_X1 port map( A1 => n897, A2 => n645, B1 => n929, B2 => n642, 
                           C1 => n865, C2 => n639, ZN => n5679);
   U2201 : OAI222_X1 port map( A1 => n1953, A2 => n483, B1 => n1985, B2 => n480
                           , C1 => n1921, C2 => n477, ZN => n5688);
   U2202 : OAI222_X1 port map( A1 => n2305, A2 => n65, B1 => n2337, B2 => n62, 
                           C1 => n2273, C2 => n59, ZN => n5697);
   U2203 : OAI222_X1 port map( A1 => n193, A2 => n1423, B1 => n225, B2 => n1420
                           , C1 => n161, C2 => n1417, ZN => n4227);
   U2204 : OAI222_X1 port map( A1 => n897, A2 => n1357, B1 => n929, B2 => n1354
                           , C1 => n865, C2 => n1351, ZN => n4236);
   U2205 : OAI222_X1 port map( A1 => n1953, A2 => n1195, B1 => n1985, B2 => 
                           n1192, C1 => n1921, C2 => n1189, ZN => n4245);
   U2206 : OAI222_X1 port map( A1 => n2305, A2 => n777, B1 => n2337, B2 => n774
                           , C1 => n2273, C2 => n771, ZN => n4254);
   U2207 : OAI222_X1 port map( A1 => n192, A2 => n711, B1 => n224, B2 => n708, 
                           C1 => n160, C2 => n705, ZN => n5629);
   U2208 : OAI222_X1 port map( A1 => n896, A2 => n645, B1 => n928, B2 => n642, 
                           C1 => n864, C2 => n639, ZN => n5638);
   U2209 : OAI222_X1 port map( A1 => n1952, A2 => n483, B1 => n1984, B2 => n480
                           , C1 => n1920, C2 => n477, ZN => n5647);
   U2210 : OAI222_X1 port map( A1 => n2304, A2 => n65, B1 => n2336, B2 => n62, 
                           C1 => n2272, C2 => n59, ZN => n5656);
   U2211 : OAI222_X1 port map( A1 => n192, A2 => n1423, B1 => n224, B2 => n1420
                           , C1 => n160, C2 => n1417, ZN => n4186);
   U2212 : OAI222_X1 port map( A1 => n896, A2 => n1357, B1 => n928, B2 => n1354
                           , C1 => n864, C2 => n1351, ZN => n4195);
   U2213 : OAI222_X1 port map( A1 => n1952, A2 => n1195, B1 => n1984, B2 => 
                           n1192, C1 => n1920, C2 => n1189, ZN => n4204);
   U2214 : OAI222_X1 port map( A1 => n2304, A2 => n777, B1 => n2336, B2 => n774
                           , C1 => n2272, C2 => n771, ZN => n4213);
   U2215 : OAI222_X1 port map( A1 => n191, A2 => n711, B1 => n223, B2 => n708, 
                           C1 => n159, C2 => n705, ZN => n5588);
   U2216 : OAI222_X1 port map( A1 => n895, A2 => n645, B1 => n927, B2 => n642, 
                           C1 => n863, C2 => n639, ZN => n5597);
   U2217 : OAI222_X1 port map( A1 => n1951, A2 => n483, B1 => n1983, B2 => n480
                           , C1 => n1919, C2 => n477, ZN => n5606);
   U2218 : OAI222_X1 port map( A1 => n2303, A2 => n65, B1 => n2335, B2 => n62, 
                           C1 => n2271, C2 => n59, ZN => n5615);
   U2219 : OAI222_X1 port map( A1 => n191, A2 => n1423, B1 => n223, B2 => n1420
                           , C1 => n159, C2 => n1417, ZN => n4145);
   U2220 : OAI222_X1 port map( A1 => n895, A2 => n1357, B1 => n927, B2 => n1354
                           , C1 => n863, C2 => n1351, ZN => n4154);
   U2221 : OAI222_X1 port map( A1 => n1951, A2 => n1195, B1 => n1983, B2 => 
                           n1192, C1 => n1919, C2 => n1189, ZN => n4163);
   U2222 : OAI222_X1 port map( A1 => n2303, A2 => n777, B1 => n2335, B2 => n774
                           , C1 => n2271, C2 => n771, ZN => n4172);
   U2223 : OAI222_X1 port map( A1 => n190, A2 => n711, B1 => n222, B2 => n708, 
                           C1 => n158, C2 => n705, ZN => n5547);
   U2224 : OAI222_X1 port map( A1 => n894, A2 => n645, B1 => n926, B2 => n642, 
                           C1 => n862, C2 => n639, ZN => n5556);
   U2225 : OAI222_X1 port map( A1 => n1950, A2 => n483, B1 => n1982, B2 => n480
                           , C1 => n1918, C2 => n477, ZN => n5565);
   U2226 : OAI222_X1 port map( A1 => n2302, A2 => n65, B1 => n2334, B2 => n62, 
                           C1 => n2270, C2 => n59, ZN => n5574);
   U2227 : OAI222_X1 port map( A1 => n190, A2 => n1423, B1 => n222, B2 => n1420
                           , C1 => n158, C2 => n1417, ZN => n4104);
   U2228 : OAI222_X1 port map( A1 => n894, A2 => n1357, B1 => n926, B2 => n1354
                           , C1 => n862, C2 => n1351, ZN => n4113);
   U2229 : OAI222_X1 port map( A1 => n1950, A2 => n1195, B1 => n1982, B2 => 
                           n1192, C1 => n1918, C2 => n1189, ZN => n4122);
   U2230 : OAI222_X1 port map( A1 => n2302, A2 => n777, B1 => n2334, B2 => n774
                           , C1 => n2270, C2 => n771, ZN => n4131);
   U2231 : OAI222_X1 port map( A1 => n189, A2 => n711, B1 => n221, B2 => n708, 
                           C1 => n157, C2 => n705, ZN => n5506);
   U2232 : OAI222_X1 port map( A1 => n893, A2 => n645, B1 => n925, B2 => n642, 
                           C1 => n861, C2 => n639, ZN => n5515);
   U2233 : OAI222_X1 port map( A1 => n1949, A2 => n483, B1 => n1981, B2 => n480
                           , C1 => n1917, C2 => n477, ZN => n5524);
   U2234 : OAI222_X1 port map( A1 => n2301, A2 => n65, B1 => n2333, B2 => n62, 
                           C1 => n2269, C2 => n59, ZN => n5533);
   U2235 : OAI222_X1 port map( A1 => n189, A2 => n1423, B1 => n221, B2 => n1420
                           , C1 => n157, C2 => n1417, ZN => n4063);
   U2236 : OAI222_X1 port map( A1 => n893, A2 => n1357, B1 => n925, B2 => n1354
                           , C1 => n861, C2 => n1351, ZN => n4072);
   U2237 : OAI222_X1 port map( A1 => n1949, A2 => n1195, B1 => n1981, B2 => 
                           n1192, C1 => n1917, C2 => n1189, ZN => n4081);
   U2238 : OAI222_X1 port map( A1 => n2301, A2 => n777, B1 => n2333, B2 => n774
                           , C1 => n2269, C2 => n771, ZN => n4090);
   U2239 : OAI222_X1 port map( A1 => n188, A2 => n711, B1 => n220, B2 => n708, 
                           C1 => n156, C2 => n705, ZN => n5465);
   U2240 : OAI222_X1 port map( A1 => n892, A2 => n645, B1 => n924, B2 => n642, 
                           C1 => n860, C2 => n639, ZN => n5474);
   U2241 : OAI222_X1 port map( A1 => n1948, A2 => n483, B1 => n1980, B2 => n480
                           , C1 => n1916, C2 => n477, ZN => n5483);
   U2242 : OAI222_X1 port map( A1 => n2300, A2 => n65, B1 => n2332, B2 => n62, 
                           C1 => n2268, C2 => n59, ZN => n5492);
   U2243 : OAI222_X1 port map( A1 => n188, A2 => n1423, B1 => n220, B2 => n1420
                           , C1 => n156, C2 => n1417, ZN => n4022);
   U2244 : OAI222_X1 port map( A1 => n892, A2 => n1357, B1 => n924, B2 => n1354
                           , C1 => n860, C2 => n1351, ZN => n4031);
   U2245 : OAI222_X1 port map( A1 => n1948, A2 => n1195, B1 => n1980, B2 => 
                           n1192, C1 => n1916, C2 => n1189, ZN => n4040);
   U2246 : OAI222_X1 port map( A1 => n2300, A2 => n777, B1 => n2332, B2 => n774
                           , C1 => n2268, C2 => n771, ZN => n4049);
   U2247 : OAI222_X1 port map( A1 => n187, A2 => n711, B1 => n219, B2 => n708, 
                           C1 => n155, C2 => n705, ZN => n5424);
   U2248 : OAI222_X1 port map( A1 => n891, A2 => n645, B1 => n923, B2 => n642, 
                           C1 => n859, C2 => n639, ZN => n5433);
   U2249 : OAI222_X1 port map( A1 => n1947, A2 => n483, B1 => n1979, B2 => n480
                           , C1 => n1915, C2 => n477, ZN => n5442);
   U2250 : OAI222_X1 port map( A1 => n2299, A2 => n65, B1 => n2331, B2 => n62, 
                           C1 => n2267, C2 => n59, ZN => n5451);
   U2251 : OAI222_X1 port map( A1 => n187, A2 => n1423, B1 => n219, B2 => n1420
                           , C1 => n155, C2 => n1417, ZN => n3981);
   U2252 : OAI222_X1 port map( A1 => n891, A2 => n1357, B1 => n923, B2 => n1354
                           , C1 => n859, C2 => n1351, ZN => n3990);
   U2253 : OAI222_X1 port map( A1 => n1947, A2 => n1195, B1 => n1979, B2 => 
                           n1192, C1 => n1915, C2 => n1189, ZN => n3999);
   U2254 : OAI222_X1 port map( A1 => n2299, A2 => n777, B1 => n2331, B2 => n774
                           , C1 => n2267, C2 => n771, ZN => n4008);
   U2255 : OAI222_X1 port map( A1 => n186, A2 => n711, B1 => n218, B2 => n708, 
                           C1 => n154, C2 => n705, ZN => n5383);
   U2256 : OAI222_X1 port map( A1 => n890, A2 => n645, B1 => n922, B2 => n642, 
                           C1 => n858, C2 => n639, ZN => n5392);
   U2257 : OAI222_X1 port map( A1 => n1946, A2 => n483, B1 => n1978, B2 => n480
                           , C1 => n1914, C2 => n477, ZN => n5401);
   U2258 : OAI222_X1 port map( A1 => n2298, A2 => n65, B1 => n2330, B2 => n62, 
                           C1 => n2266, C2 => n59, ZN => n5410);
   U2259 : OAI222_X1 port map( A1 => n186, A2 => n1423, B1 => n218, B2 => n1420
                           , C1 => n154, C2 => n1417, ZN => n3940);
   U2260 : OAI222_X1 port map( A1 => n890, A2 => n1357, B1 => n922, B2 => n1354
                           , C1 => n858, C2 => n1351, ZN => n3949);
   U2261 : OAI222_X1 port map( A1 => n1946, A2 => n1195, B1 => n1978, B2 => 
                           n1192, C1 => n1914, C2 => n1189, ZN => n3958);
   U2262 : OAI222_X1 port map( A1 => n2298, A2 => n777, B1 => n2330, B2 => n774
                           , C1 => n2266, C2 => n771, ZN => n3967);
   U2263 : OAI222_X1 port map( A1 => n185, A2 => n711, B1 => n217, B2 => n708, 
                           C1 => n153, C2 => n705, ZN => n5342);
   U2264 : OAI222_X1 port map( A1 => n889, A2 => n645, B1 => n921, B2 => n642, 
                           C1 => n857, C2 => n639, ZN => n5351);
   U2265 : OAI222_X1 port map( A1 => n1945, A2 => n483, B1 => n1977, B2 => n480
                           , C1 => n1913, C2 => n477, ZN => n5360);
   U2266 : OAI222_X1 port map( A1 => n2297, A2 => n65, B1 => n2329, B2 => n62, 
                           C1 => n2265, C2 => n59, ZN => n5369);
   U2267 : OAI222_X1 port map( A1 => n185, A2 => n1423, B1 => n217, B2 => n1420
                           , C1 => n153, C2 => n1417, ZN => n3899);
   U2268 : OAI222_X1 port map( A1 => n889, A2 => n1357, B1 => n921, B2 => n1354
                           , C1 => n857, C2 => n1351, ZN => n3908);
   U2269 : OAI222_X1 port map( A1 => n1945, A2 => n1195, B1 => n1977, B2 => 
                           n1192, C1 => n1913, C2 => n1189, ZN => n3917);
   U2270 : OAI222_X1 port map( A1 => n2297, A2 => n777, B1 => n2329, B2 => n774
                           , C1 => n2265, C2 => n771, ZN => n3926);
   U2271 : OAI222_X1 port map( A1 => n184, A2 => n711, B1 => n216, B2 => n708, 
                           C1 => n152, C2 => n705, ZN => n5301);
   U2272 : OAI222_X1 port map( A1 => n888, A2 => n645, B1 => n920, B2 => n642, 
                           C1 => n856, C2 => n639, ZN => n5310);
   U2273 : OAI222_X1 port map( A1 => n1944, A2 => n483, B1 => n1976, B2 => n480
                           , C1 => n1912, C2 => n477, ZN => n5319);
   U2274 : OAI222_X1 port map( A1 => n2296, A2 => n65, B1 => n2328, B2 => n62, 
                           C1 => n2264, C2 => n59, ZN => n5328);
   U2275 : OAI222_X1 port map( A1 => n184, A2 => n1423, B1 => n216, B2 => n1420
                           , C1 => n152, C2 => n1417, ZN => n3858);
   U2276 : OAI222_X1 port map( A1 => n888, A2 => n1357, B1 => n920, B2 => n1354
                           , C1 => n856, C2 => n1351, ZN => n3867);
   U2277 : OAI222_X1 port map( A1 => n1944, A2 => n1195, B1 => n1976, B2 => 
                           n1192, C1 => n1912, C2 => n1189, ZN => n3876);
   U2278 : OAI222_X1 port map( A1 => n2296, A2 => n777, B1 => n2328, B2 => n774
                           , C1 => n2264, C2 => n771, ZN => n3885);
   U2279 : OAI222_X1 port map( A1 => n183, A2 => n712, B1 => n215, B2 => n709, 
                           C1 => n151, C2 => n706, ZN => n5260);
   U2280 : OAI222_X1 port map( A1 => n887, A2 => n646, B1 => n919, B2 => n643, 
                           C1 => n855, C2 => n640, ZN => n5269);
   U2281 : OAI222_X1 port map( A1 => n1943, A2 => n484, B1 => n1975, B2 => n481
                           , C1 => n1911, C2 => n478, ZN => n5278);
   U2282 : OAI222_X1 port map( A1 => n2295, A2 => n66, B1 => n2327, B2 => n63, 
                           C1 => n2263, C2 => n60, ZN => n5287);
   U2283 : OAI222_X1 port map( A1 => n183, A2 => n1424, B1 => n215, B2 => n1421
                           , C1 => n151, C2 => n1418, ZN => n3817);
   U2284 : OAI222_X1 port map( A1 => n887, A2 => n1358, B1 => n919, B2 => n1355
                           , C1 => n855, C2 => n1352, ZN => n3826);
   U2285 : OAI222_X1 port map( A1 => n1943, A2 => n1196, B1 => n1975, B2 => 
                           n1193, C1 => n1911, C2 => n1190, ZN => n3835);
   U2286 : OAI222_X1 port map( A1 => n2295, A2 => n778, B1 => n2327, B2 => n775
                           , C1 => n2263, C2 => n772, ZN => n3844);
   U2287 : OAI222_X1 port map( A1 => n182, A2 => n712, B1 => n214, B2 => n709, 
                           C1 => n150, C2 => n706, ZN => n5219);
   U2288 : OAI222_X1 port map( A1 => n886, A2 => n646, B1 => n918, B2 => n643, 
                           C1 => n854, C2 => n640, ZN => n5228);
   U2289 : OAI222_X1 port map( A1 => n1942, A2 => n484, B1 => n1974, B2 => n481
                           , C1 => n1910, C2 => n478, ZN => n5237);
   U2290 : OAI222_X1 port map( A1 => n2294, A2 => n66, B1 => n2326, B2 => n63, 
                           C1 => n2262, C2 => n60, ZN => n5246);
   U2291 : OAI222_X1 port map( A1 => n182, A2 => n1424, B1 => n214, B2 => n1421
                           , C1 => n150, C2 => n1418, ZN => n3776);
   U2292 : OAI222_X1 port map( A1 => n886, A2 => n1358, B1 => n918, B2 => n1355
                           , C1 => n854, C2 => n1352, ZN => n3785);
   U2293 : OAI222_X1 port map( A1 => n1942, A2 => n1196, B1 => n1974, B2 => 
                           n1193, C1 => n1910, C2 => n1190, ZN => n3794);
   U2294 : OAI222_X1 port map( A1 => n2294, A2 => n778, B1 => n2326, B2 => n775
                           , C1 => n2262, C2 => n772, ZN => n3803);
   U2295 : OAI222_X1 port map( A1 => n181, A2 => n712, B1 => n213, B2 => n709, 
                           C1 => n149, C2 => n706, ZN => n5178);
   U2296 : OAI222_X1 port map( A1 => n885, A2 => n646, B1 => n917, B2 => n643, 
                           C1 => n853, C2 => n640, ZN => n5187);
   U2297 : OAI222_X1 port map( A1 => n1941, A2 => n484, B1 => n1973, B2 => n481
                           , C1 => n1909, C2 => n478, ZN => n5196);
   U2298 : OAI222_X1 port map( A1 => n2293, A2 => n66, B1 => n2325, B2 => n63, 
                           C1 => n2261, C2 => n60, ZN => n5205);
   U2299 : OAI222_X1 port map( A1 => n181, A2 => n1424, B1 => n213, B2 => n1421
                           , C1 => n149, C2 => n1418, ZN => n3735);
   U2300 : OAI222_X1 port map( A1 => n885, A2 => n1358, B1 => n917, B2 => n1355
                           , C1 => n853, C2 => n1352, ZN => n3744);
   U2301 : OAI222_X1 port map( A1 => n1941, A2 => n1196, B1 => n1973, B2 => 
                           n1193, C1 => n1909, C2 => n1190, ZN => n3753);
   U2302 : OAI222_X1 port map( A1 => n2293, A2 => n778, B1 => n2325, B2 => n775
                           , C1 => n2261, C2 => n772, ZN => n3762);
   U2303 : OAI222_X1 port map( A1 => n180, A2 => n712, B1 => n212, B2 => n709, 
                           C1 => n148, C2 => n706, ZN => n5137);
   U2304 : OAI222_X1 port map( A1 => n884, A2 => n646, B1 => n916, B2 => n643, 
                           C1 => n852, C2 => n640, ZN => n5146);
   U2305 : OAI222_X1 port map( A1 => n1940, A2 => n484, B1 => n1972, B2 => n481
                           , C1 => n1908, C2 => n478, ZN => n5155);
   U2306 : OAI222_X1 port map( A1 => n2292, A2 => n66, B1 => n2324, B2 => n63, 
                           C1 => n2260, C2 => n60, ZN => n5164);
   U2307 : OAI222_X1 port map( A1 => n180, A2 => n1424, B1 => n212, B2 => n1421
                           , C1 => n148, C2 => n1418, ZN => n3694);
   U2308 : OAI222_X1 port map( A1 => n884, A2 => n1358, B1 => n916, B2 => n1355
                           , C1 => n852, C2 => n1352, ZN => n3703);
   U2309 : OAI222_X1 port map( A1 => n1940, A2 => n1196, B1 => n1972, B2 => 
                           n1193, C1 => n1908, C2 => n1190, ZN => n3712);
   U2310 : OAI222_X1 port map( A1 => n2292, A2 => n778, B1 => n2324, B2 => n775
                           , C1 => n2260, C2 => n772, ZN => n3721);
   U2311 : OAI222_X1 port map( A1 => n179, A2 => n712, B1 => n211, B2 => n709, 
                           C1 => n147, C2 => n706, ZN => n5096);
   U2312 : OAI222_X1 port map( A1 => n883, A2 => n646, B1 => n915, B2 => n643, 
                           C1 => n851, C2 => n640, ZN => n5105);
   U2313 : OAI222_X1 port map( A1 => n1939, A2 => n484, B1 => n1971, B2 => n481
                           , C1 => n1907, C2 => n478, ZN => n5114);
   U2314 : OAI222_X1 port map( A1 => n2291, A2 => n66, B1 => n2323, B2 => n63, 
                           C1 => n2259, C2 => n60, ZN => n5123);
   U2315 : OAI222_X1 port map( A1 => n179, A2 => n1424, B1 => n211, B2 => n1421
                           , C1 => n147, C2 => n1418, ZN => n3653);
   U2316 : OAI222_X1 port map( A1 => n883, A2 => n1358, B1 => n915, B2 => n1355
                           , C1 => n851, C2 => n1352, ZN => n3662);
   U2317 : OAI222_X1 port map( A1 => n1939, A2 => n1196, B1 => n1971, B2 => 
                           n1193, C1 => n1907, C2 => n1190, ZN => n3671);
   U2318 : OAI222_X1 port map( A1 => n2291, A2 => n778, B1 => n2323, B2 => n775
                           , C1 => n2259, C2 => n772, ZN => n3680);
   U2319 : OAI222_X1 port map( A1 => n178, A2 => n712, B1 => n210, B2 => n709, 
                           C1 => n146, C2 => n706, ZN => n5055);
   U2320 : OAI222_X1 port map( A1 => n882, A2 => n646, B1 => n914, B2 => n643, 
                           C1 => n850, C2 => n640, ZN => n5064);
   U2321 : OAI222_X1 port map( A1 => n1938, A2 => n484, B1 => n1970, B2 => n481
                           , C1 => n1906, C2 => n478, ZN => n5073);
   U2322 : OAI222_X1 port map( A1 => n2290, A2 => n66, B1 => n2322, B2 => n63, 
                           C1 => n2258, C2 => n60, ZN => n5082);
   U2323 : OAI222_X1 port map( A1 => n178, A2 => n1424, B1 => n210, B2 => n1421
                           , C1 => n146, C2 => n1418, ZN => n3612);
   U2324 : OAI222_X1 port map( A1 => n882, A2 => n1358, B1 => n914, B2 => n1355
                           , C1 => n850, C2 => n1352, ZN => n3621);
   U2325 : OAI222_X1 port map( A1 => n1938, A2 => n1196, B1 => n1970, B2 => 
                           n1193, C1 => n1906, C2 => n1190, ZN => n3630);
   U2326 : OAI222_X1 port map( A1 => n2290, A2 => n778, B1 => n2322, B2 => n775
                           , C1 => n2258, C2 => n772, ZN => n3639);
   U2327 : OAI222_X1 port map( A1 => n177, A2 => n712, B1 => n209, B2 => n709, 
                           C1 => n145, C2 => n706, ZN => n5014);
   U2328 : OAI222_X1 port map( A1 => n881, A2 => n646, B1 => n913, B2 => n643, 
                           C1 => n849, C2 => n640, ZN => n5023);
   U2329 : OAI222_X1 port map( A1 => n1937, A2 => n484, B1 => n1969, B2 => n481
                           , C1 => n1905, C2 => n478, ZN => n5032);
   U2330 : OAI222_X1 port map( A1 => n2289, A2 => n66, B1 => n2321, B2 => n63, 
                           C1 => n2257, C2 => n60, ZN => n5041);
   U2331 : OAI222_X1 port map( A1 => n177, A2 => n1424, B1 => n209, B2 => n1421
                           , C1 => n145, C2 => n1418, ZN => n3571);
   U2332 : OAI222_X1 port map( A1 => n881, A2 => n1358, B1 => n913, B2 => n1355
                           , C1 => n849, C2 => n1352, ZN => n3580);
   U2333 : OAI222_X1 port map( A1 => n1937, A2 => n1196, B1 => n1969, B2 => 
                           n1193, C1 => n1905, C2 => n1190, ZN => n3589);
   U2334 : OAI222_X1 port map( A1 => n2289, A2 => n778, B1 => n2321, B2 => n775
                           , C1 => n2257, C2 => n772, ZN => n3598);
   U2335 : OAI222_X1 port map( A1 => n176, A2 => n712, B1 => n208, B2 => n709, 
                           C1 => n144, C2 => n706, ZN => n4885);
   U2336 : OAI222_X1 port map( A1 => n880, A2 => n646, B1 => n912, B2 => n643, 
                           C1 => n848, C2 => n640, ZN => n4916);
   U2337 : OAI222_X1 port map( A1 => n1936, A2 => n484, B1 => n1968, B2 => n481
                           , C1 => n1904, C2 => n478, ZN => n4947);
   U2338 : OAI222_X1 port map( A1 => n2288, A2 => n66, B1 => n2320, B2 => n63, 
                           C1 => n2256, C2 => n60, ZN => n4978);
   U2339 : OAI222_X1 port map( A1 => n176, A2 => n1424, B1 => n208, B2 => n1421
                           , C1 => n144, C2 => n1418, ZN => n3442);
   U2340 : OAI222_X1 port map( A1 => n880, A2 => n1358, B1 => n912, B2 => n1355
                           , C1 => n848, C2 => n1352, ZN => n3473);
   U2341 : OAI222_X1 port map( A1 => n1936, A2 => n1196, B1 => n1968, B2 => 
                           n1193, C1 => n1904, C2 => n1190, ZN => n3504);
   U2342 : OAI222_X1 port map( A1 => n2288, A2 => n778, B1 => n2320, B2 => n775
                           , C1 => n2256, C2 => n772, ZN => n3535);
   U2343 : OAI222_X1 port map( A1 => n559, A2 => n677, B1 => n591, B2 => n674, 
                           C1 => n527, C2 => n671, ZN => n6258);
   U2344 : OAI222_X1 port map( A1 => n1263, A2 => n611, B1 => n1295, B2 => n608
                           , C1 => n1231, C2 => n605, ZN => n6282);
   U2345 : OAI222_X1 port map( A1 => n559, A2 => n1389, B1 => n591, B2 => n1386
                           , C1 => n527, C2 => n1383, ZN => n4815);
   U2346 : OAI222_X1 port map( A1 => n1263, A2 => n1323, B1 => n1295, B2 => 
                           n1320, C1 => n1231, C2 => n1317, ZN => n4839);
   U2347 : OAI222_X1 port map( A1 => n558, A2 => n677, B1 => n590, B2 => n674, 
                           C1 => n526, C2 => n671, ZN => n6205);
   U2348 : OAI222_X1 port map( A1 => n1262, A2 => n611, B1 => n1294, B2 => n608
                           , C1 => n1230, C2 => n605, ZN => n6214);
   U2349 : OAI222_X1 port map( A1 => n558, A2 => n1389, B1 => n590, B2 => n1386
                           , C1 => n526, C2 => n1383, ZN => n4762);
   U2350 : OAI222_X1 port map( A1 => n1262, A2 => n1323, B1 => n1294, B2 => 
                           n1320, C1 => n1230, C2 => n1317, ZN => n4771);
   U2351 : OAI222_X1 port map( A1 => n557, A2 => n677, B1 => n589, B2 => n674, 
                           C1 => n525, C2 => n671, ZN => n6164);
   U2352 : OAI222_X1 port map( A1 => n1261, A2 => n611, B1 => n1293, B2 => n608
                           , C1 => n1229, C2 => n605, ZN => n6173);
   U2353 : OAI222_X1 port map( A1 => n557, A2 => n1389, B1 => n589, B2 => n1386
                           , C1 => n525, C2 => n1383, ZN => n4721);
   U2354 : OAI222_X1 port map( A1 => n1261, A2 => n1323, B1 => n1293, B2 => 
                           n1320, C1 => n1229, C2 => n1317, ZN => n4730);
   U2355 : OAI222_X1 port map( A1 => n556, A2 => n677, B1 => n588, B2 => n674, 
                           C1 => n524, C2 => n671, ZN => n6123);
   U2356 : OAI222_X1 port map( A1 => n1260, A2 => n611, B1 => n1292, B2 => n608
                           , C1 => n1228, C2 => n605, ZN => n6132);
   U2357 : OAI222_X1 port map( A1 => n556, A2 => n1389, B1 => n588, B2 => n1386
                           , C1 => n524, C2 => n1383, ZN => n4680);
   U2358 : OAI222_X1 port map( A1 => n1260, A2 => n1323, B1 => n1292, B2 => 
                           n1320, C1 => n1228, C2 => n1317, ZN => n4689);
   U2359 : OAI222_X1 port map( A1 => n555, A2 => n677, B1 => n587, B2 => n674, 
                           C1 => n523, C2 => n671, ZN => n6082);
   U2360 : OAI222_X1 port map( A1 => n1259, A2 => n611, B1 => n1291, B2 => n608
                           , C1 => n1227, C2 => n605, ZN => n6091);
   U2361 : OAI222_X1 port map( A1 => n555, A2 => n1389, B1 => n587, B2 => n1386
                           , C1 => n523, C2 => n1383, ZN => n4639);
   U2362 : OAI222_X1 port map( A1 => n1259, A2 => n1323, B1 => n1291, B2 => 
                           n1320, C1 => n1227, C2 => n1317, ZN => n4648);
   U2363 : OAI222_X1 port map( A1 => n554, A2 => n677, B1 => n586, B2 => n674, 
                           C1 => n522, C2 => n671, ZN => n6041);
   U2364 : OAI222_X1 port map( A1 => n1258, A2 => n611, B1 => n1290, B2 => n608
                           , C1 => n1226, C2 => n605, ZN => n6050);
   U2365 : OAI222_X1 port map( A1 => n554, A2 => n1389, B1 => n586, B2 => n1386
                           , C1 => n522, C2 => n1383, ZN => n4598);
   U2366 : OAI222_X1 port map( A1 => n1258, A2 => n1323, B1 => n1290, B2 => 
                           n1320, C1 => n1226, C2 => n1317, ZN => n4607);
   U2367 : OAI222_X1 port map( A1 => n553, A2 => n677, B1 => n585, B2 => n674, 
                           C1 => n521, C2 => n671, ZN => n6000);
   U2368 : OAI222_X1 port map( A1 => n1257, A2 => n611, B1 => n1289, B2 => n608
                           , C1 => n1225, C2 => n605, ZN => n6009);
   U2369 : OAI222_X1 port map( A1 => n553, A2 => n1389, B1 => n585, B2 => n1386
                           , C1 => n521, C2 => n1383, ZN => n4557);
   U2370 : OAI222_X1 port map( A1 => n1257, A2 => n1323, B1 => n1289, B2 => 
                           n1320, C1 => n1225, C2 => n1317, ZN => n4566);
   U2371 : OAI222_X1 port map( A1 => n552, A2 => n677, B1 => n584, B2 => n674, 
                           C1 => n520, C2 => n671, ZN => n5959);
   U2372 : OAI222_X1 port map( A1 => n1256, A2 => n611, B1 => n1288, B2 => n608
                           , C1 => n1224, C2 => n605, ZN => n5968);
   U2373 : OAI222_X1 port map( A1 => n552, A2 => n1389, B1 => n584, B2 => n1386
                           , C1 => n520, C2 => n1383, ZN => n4516);
   U2374 : OAI222_X1 port map( A1 => n1256, A2 => n1323, B1 => n1288, B2 => 
                           n1320, C1 => n1224, C2 => n1317, ZN => n4525);
   U2375 : OAI222_X1 port map( A1 => n551, A2 => n677, B1 => n583, B2 => n674, 
                           C1 => n519, C2 => n671, ZN => n5918);
   U2376 : OAI222_X1 port map( A1 => n1255, A2 => n611, B1 => n1287, B2 => n608
                           , C1 => n1223, C2 => n605, ZN => n5927);
   U2377 : OAI222_X1 port map( A1 => n551, A2 => n1389, B1 => n583, B2 => n1386
                           , C1 => n519, C2 => n1383, ZN => n4475);
   U2378 : OAI222_X1 port map( A1 => n1255, A2 => n1323, B1 => n1287, B2 => 
                           n1320, C1 => n1223, C2 => n1317, ZN => n4484);
   U2379 : OAI222_X1 port map( A1 => n550, A2 => n677, B1 => n582, B2 => n674, 
                           C1 => n518, C2 => n671, ZN => n5877);
   U2380 : OAI222_X1 port map( A1 => n1254, A2 => n611, B1 => n1286, B2 => n608
                           , C1 => n1222, C2 => n605, ZN => n5886);
   U2381 : OAI222_X1 port map( A1 => n550, A2 => n1389, B1 => n582, B2 => n1386
                           , C1 => n518, C2 => n1383, ZN => n4434);
   U2382 : OAI222_X1 port map( A1 => n1254, A2 => n1323, B1 => n1286, B2 => 
                           n1320, C1 => n1222, C2 => n1317, ZN => n4443);
   U2383 : OAI222_X1 port map( A1 => n549, A2 => n677, B1 => n581, B2 => n674, 
                           C1 => n517, C2 => n671, ZN => n5836);
   U2384 : OAI222_X1 port map( A1 => n1253, A2 => n611, B1 => n1285, B2 => n608
                           , C1 => n1221, C2 => n605, ZN => n5845);
   U2385 : OAI222_X1 port map( A1 => n549, A2 => n1389, B1 => n581, B2 => n1386
                           , C1 => n517, C2 => n1383, ZN => n4393);
   U2386 : OAI222_X1 port map( A1 => n1253, A2 => n1323, B1 => n1285, B2 => 
                           n1320, C1 => n1221, C2 => n1317, ZN => n4402);
   U2387 : OAI222_X1 port map( A1 => n548, A2 => n677, B1 => n580, B2 => n674, 
                           C1 => n516, C2 => n671, ZN => n5795);
   U2388 : OAI222_X1 port map( A1 => n1252, A2 => n611, B1 => n1284, B2 => n608
                           , C1 => n1220, C2 => n605, ZN => n5804);
   U2389 : OAI222_X1 port map( A1 => n548, A2 => n1389, B1 => n580, B2 => n1386
                           , C1 => n516, C2 => n1383, ZN => n4352);
   U2390 : OAI222_X1 port map( A1 => n1252, A2 => n1323, B1 => n1284, B2 => 
                           n1320, C1 => n1220, C2 => n1317, ZN => n4361);
   U2391 : OAI222_X1 port map( A1 => n547, A2 => n678, B1 => n579, B2 => n675, 
                           C1 => n515, C2 => n672, ZN => n5754);
   U2392 : OAI222_X1 port map( A1 => n1251, A2 => n612, B1 => n1283, B2 => n609
                           , C1 => n1219, C2 => n606, ZN => n5763);
   U2393 : OAI222_X1 port map( A1 => n547, A2 => n1390, B1 => n579, B2 => n1387
                           , C1 => n515, C2 => n1384, ZN => n4311);
   U2394 : OAI222_X1 port map( A1 => n1251, A2 => n1324, B1 => n1283, B2 => 
                           n1321, C1 => n1219, C2 => n1318, ZN => n4320);
   U2395 : OAI222_X1 port map( A1 => n546, A2 => n678, B1 => n578, B2 => n675, 
                           C1 => n514, C2 => n672, ZN => n5713);
   U2396 : OAI222_X1 port map( A1 => n1250, A2 => n612, B1 => n1282, B2 => n609
                           , C1 => n1218, C2 => n606, ZN => n5722);
   U2397 : OAI222_X1 port map( A1 => n546, A2 => n1390, B1 => n578, B2 => n1387
                           , C1 => n514, C2 => n1384, ZN => n4270);
   U2398 : OAI222_X1 port map( A1 => n1250, A2 => n1324, B1 => n1282, B2 => 
                           n1321, C1 => n1218, C2 => n1318, ZN => n4279);
   U2399 : OAI222_X1 port map( A1 => n545, A2 => n678, B1 => n577, B2 => n675, 
                           C1 => n513, C2 => n672, ZN => n5672);
   U2400 : OAI222_X1 port map( A1 => n1249, A2 => n612, B1 => n1281, B2 => n609
                           , C1 => n1217, C2 => n606, ZN => n5681);
   U2401 : OAI222_X1 port map( A1 => n545, A2 => n1390, B1 => n577, B2 => n1387
                           , C1 => n513, C2 => n1384, ZN => n4229);
   U2402 : OAI222_X1 port map( A1 => n1249, A2 => n1324, B1 => n1281, B2 => 
                           n1321, C1 => n1217, C2 => n1318, ZN => n4238);
   U2403 : OAI222_X1 port map( A1 => n544, A2 => n678, B1 => n576, B2 => n675, 
                           C1 => n512, C2 => n672, ZN => n5631);
   U2404 : OAI222_X1 port map( A1 => n1248, A2 => n612, B1 => n1280, B2 => n609
                           , C1 => n1216, C2 => n606, ZN => n5640);
   U2405 : OAI222_X1 port map( A1 => n544, A2 => n1390, B1 => n576, B2 => n1387
                           , C1 => n512, C2 => n1384, ZN => n4188);
   U2406 : OAI222_X1 port map( A1 => n1248, A2 => n1324, B1 => n1280, B2 => 
                           n1321, C1 => n1216, C2 => n1318, ZN => n4197);
   U2407 : OAI222_X1 port map( A1 => n543, A2 => n678, B1 => n575, B2 => n675, 
                           C1 => n511, C2 => n672, ZN => n5590);
   U2408 : OAI222_X1 port map( A1 => n1247, A2 => n612, B1 => n1279, B2 => n609
                           , C1 => n1215, C2 => n606, ZN => n5599);
   U2409 : OAI222_X1 port map( A1 => n543, A2 => n1390, B1 => n575, B2 => n1387
                           , C1 => n511, C2 => n1384, ZN => n4147);
   U2410 : OAI222_X1 port map( A1 => n1247, A2 => n1324, B1 => n1279, B2 => 
                           n1321, C1 => n1215, C2 => n1318, ZN => n4156);
   U2411 : OAI222_X1 port map( A1 => n542, A2 => n678, B1 => n574, B2 => n675, 
                           C1 => n510, C2 => n672, ZN => n5549);
   U2412 : OAI222_X1 port map( A1 => n1246, A2 => n612, B1 => n1278, B2 => n609
                           , C1 => n1214, C2 => n606, ZN => n5558);
   U2413 : OAI222_X1 port map( A1 => n542, A2 => n1390, B1 => n574, B2 => n1387
                           , C1 => n510, C2 => n1384, ZN => n4106);
   U2414 : OAI222_X1 port map( A1 => n1246, A2 => n1324, B1 => n1278, B2 => 
                           n1321, C1 => n1214, C2 => n1318, ZN => n4115);
   U2415 : OAI222_X1 port map( A1 => n541, A2 => n678, B1 => n573, B2 => n675, 
                           C1 => n509, C2 => n672, ZN => n5508);
   U2416 : OAI222_X1 port map( A1 => n1245, A2 => n612, B1 => n1277, B2 => n609
                           , C1 => n1213, C2 => n606, ZN => n5517);
   U2417 : OAI222_X1 port map( A1 => n541, A2 => n1390, B1 => n573, B2 => n1387
                           , C1 => n509, C2 => n1384, ZN => n4065);
   U2418 : OAI222_X1 port map( A1 => n1245, A2 => n1324, B1 => n1277, B2 => 
                           n1321, C1 => n1213, C2 => n1318, ZN => n4074);
   U2419 : OAI222_X1 port map( A1 => n540, A2 => n678, B1 => n572, B2 => n675, 
                           C1 => n508, C2 => n672, ZN => n5467);
   U2420 : OAI222_X1 port map( A1 => n1244, A2 => n612, B1 => n1276, B2 => n609
                           , C1 => n1212, C2 => n606, ZN => n5476);
   U2421 : OAI222_X1 port map( A1 => n540, A2 => n1390, B1 => n572, B2 => n1387
                           , C1 => n508, C2 => n1384, ZN => n4024);
   U2422 : OAI222_X1 port map( A1 => n1244, A2 => n1324, B1 => n1276, B2 => 
                           n1321, C1 => n1212, C2 => n1318, ZN => n4033);
   U2423 : OAI222_X1 port map( A1 => n539, A2 => n678, B1 => n571, B2 => n675, 
                           C1 => n507, C2 => n672, ZN => n5426);
   U2424 : OAI222_X1 port map( A1 => n1243, A2 => n612, B1 => n1275, B2 => n609
                           , C1 => n1211, C2 => n606, ZN => n5435);
   U2425 : OAI222_X1 port map( A1 => n539, A2 => n1390, B1 => n571, B2 => n1387
                           , C1 => n507, C2 => n1384, ZN => n3983);
   U2426 : OAI222_X1 port map( A1 => n1243, A2 => n1324, B1 => n1275, B2 => 
                           n1321, C1 => n1211, C2 => n1318, ZN => n3992);
   U2427 : OAI222_X1 port map( A1 => n538, A2 => n678, B1 => n570, B2 => n675, 
                           C1 => n506, C2 => n672, ZN => n5385);
   U2428 : OAI222_X1 port map( A1 => n1242, A2 => n612, B1 => n1274, B2 => n609
                           , C1 => n1210, C2 => n606, ZN => n5394);
   U2429 : OAI222_X1 port map( A1 => n538, A2 => n1390, B1 => n570, B2 => n1387
                           , C1 => n506, C2 => n1384, ZN => n3942);
   U2430 : OAI222_X1 port map( A1 => n1242, A2 => n1324, B1 => n1274, B2 => 
                           n1321, C1 => n1210, C2 => n1318, ZN => n3951);
   U2431 : OAI222_X1 port map( A1 => n537, A2 => n678, B1 => n569, B2 => n675, 
                           C1 => n505, C2 => n672, ZN => n5344);
   U2432 : OAI222_X1 port map( A1 => n1241, A2 => n612, B1 => n1273, B2 => n609
                           , C1 => n1209, C2 => n606, ZN => n5353);
   U2433 : OAI222_X1 port map( A1 => n537, A2 => n1390, B1 => n569, B2 => n1387
                           , C1 => n505, C2 => n1384, ZN => n3901);
   U2434 : OAI222_X1 port map( A1 => n1241, A2 => n1324, B1 => n1273, B2 => 
                           n1321, C1 => n1209, C2 => n1318, ZN => n3910);
   U2435 : OAI222_X1 port map( A1 => n536, A2 => n678, B1 => n568, B2 => n675, 
                           C1 => n504, C2 => n672, ZN => n5303);
   U2436 : OAI222_X1 port map( A1 => n1240, A2 => n612, B1 => n1272, B2 => n609
                           , C1 => n1208, C2 => n606, ZN => n5312);
   U2437 : OAI222_X1 port map( A1 => n536, A2 => n1390, B1 => n568, B2 => n1387
                           , C1 => n504, C2 => n1384, ZN => n3860);
   U2438 : OAI222_X1 port map( A1 => n1240, A2 => n1324, B1 => n1272, B2 => 
                           n1321, C1 => n1208, C2 => n1318, ZN => n3869);
   U2439 : OAI222_X1 port map( A1 => n535, A2 => n679, B1 => n567, B2 => n676, 
                           C1 => n503, C2 => n673, ZN => n5262);
   U2440 : OAI222_X1 port map( A1 => n1239, A2 => n613, B1 => n1271, B2 => n610
                           , C1 => n1207, C2 => n607, ZN => n5271);
   U2441 : OAI222_X1 port map( A1 => n535, A2 => n1391, B1 => n567, B2 => n1388
                           , C1 => n503, C2 => n1385, ZN => n3819);
   U2442 : OAI222_X1 port map( A1 => n1239, A2 => n1325, B1 => n1271, B2 => 
                           n1322, C1 => n1207, C2 => n1319, ZN => n3828);
   U2443 : OAI222_X1 port map( A1 => n534, A2 => n679, B1 => n566, B2 => n676, 
                           C1 => n502, C2 => n673, ZN => n5221);
   U2444 : OAI222_X1 port map( A1 => n1238, A2 => n613, B1 => n1270, B2 => n610
                           , C1 => n1206, C2 => n607, ZN => n5230);
   U2445 : OAI222_X1 port map( A1 => n534, A2 => n1391, B1 => n566, B2 => n1388
                           , C1 => n502, C2 => n1385, ZN => n3778);
   U2446 : OAI222_X1 port map( A1 => n1238, A2 => n1325, B1 => n1270, B2 => 
                           n1322, C1 => n1206, C2 => n1319, ZN => n3787);
   U2447 : OAI222_X1 port map( A1 => n533, A2 => n679, B1 => n565, B2 => n676, 
                           C1 => n501, C2 => n673, ZN => n5180);
   U2448 : OAI222_X1 port map( A1 => n1237, A2 => n613, B1 => n1269, B2 => n610
                           , C1 => n1205, C2 => n607, ZN => n5189);
   U2449 : OAI222_X1 port map( A1 => n533, A2 => n1391, B1 => n565, B2 => n1388
                           , C1 => n501, C2 => n1385, ZN => n3737);
   U2450 : OAI222_X1 port map( A1 => n1237, A2 => n1325, B1 => n1269, B2 => 
                           n1322, C1 => n1205, C2 => n1319, ZN => n3746);
   U2451 : OAI222_X1 port map( A1 => n532, A2 => n679, B1 => n564, B2 => n676, 
                           C1 => n500, C2 => n673, ZN => n5139);
   U2452 : OAI222_X1 port map( A1 => n1236, A2 => n613, B1 => n1268, B2 => n610
                           , C1 => n1204, C2 => n607, ZN => n5148);
   U2453 : OAI222_X1 port map( A1 => n532, A2 => n1391, B1 => n564, B2 => n1388
                           , C1 => n500, C2 => n1385, ZN => n3696);
   U2454 : OAI222_X1 port map( A1 => n1236, A2 => n1325, B1 => n1268, B2 => 
                           n1322, C1 => n1204, C2 => n1319, ZN => n3705);
   U2455 : OAI222_X1 port map( A1 => n531, A2 => n679, B1 => n563, B2 => n676, 
                           C1 => n499, C2 => n673, ZN => n5098);
   U2456 : OAI222_X1 port map( A1 => n1235, A2 => n613, B1 => n1267, B2 => n610
                           , C1 => n1203, C2 => n607, ZN => n5107);
   U2457 : OAI222_X1 port map( A1 => n531, A2 => n1391, B1 => n563, B2 => n1388
                           , C1 => n499, C2 => n1385, ZN => n3655);
   U2458 : OAI222_X1 port map( A1 => n1235, A2 => n1325, B1 => n1267, B2 => 
                           n1322, C1 => n1203, C2 => n1319, ZN => n3664);
   U2459 : OAI222_X1 port map( A1 => n530, A2 => n679, B1 => n562, B2 => n676, 
                           C1 => n498, C2 => n673, ZN => n5057);
   U2460 : OAI222_X1 port map( A1 => n1234, A2 => n613, B1 => n1266, B2 => n610
                           , C1 => n1202, C2 => n607, ZN => n5066);
   U2461 : OAI222_X1 port map( A1 => n530, A2 => n1391, B1 => n562, B2 => n1388
                           , C1 => n498, C2 => n1385, ZN => n3614);
   U2462 : OAI222_X1 port map( A1 => n1234, A2 => n1325, B1 => n1266, B2 => 
                           n1322, C1 => n1202, C2 => n1319, ZN => n3623);
   U2463 : OAI222_X1 port map( A1 => n529, A2 => n679, B1 => n561, B2 => n676, 
                           C1 => n497, C2 => n673, ZN => n5016);
   U2464 : OAI222_X1 port map( A1 => n1233, A2 => n613, B1 => n1265, B2 => n610
                           , C1 => n1201, C2 => n607, ZN => n5025);
   U2465 : OAI222_X1 port map( A1 => n529, A2 => n1391, B1 => n561, B2 => n1388
                           , C1 => n497, C2 => n1385, ZN => n3573);
   U2466 : OAI222_X1 port map( A1 => n1233, A2 => n1325, B1 => n1265, B2 => 
                           n1322, C1 => n1201, C2 => n1319, ZN => n3582);
   U2467 : OAI222_X1 port map( A1 => n528, A2 => n679, B1 => n560, B2 => n676, 
                           C1 => n496, C2 => n673, ZN => n4900);
   U2468 : OAI222_X1 port map( A1 => n1232, A2 => n613, B1 => n1264, B2 => n610
                           , C1 => n1200, C2 => n607, ZN => n4931);
   U2469 : OAI222_X1 port map( A1 => n528, A2 => n1391, B1 => n560, B2 => n1388
                           , C1 => n496, C2 => n1385, ZN => n3457);
   U2470 : OAI222_X1 port map( A1 => n1232, A2 => n1325, B1 => n1264, B2 => 
                           n1322, C1 => n1200, C2 => n1319, ZN => n3488);
   U2471 : OAI222_X1 port map( A1 => n303, A2 => n701, B1 => n335, B2 => n698, 
                           C1 => n271, C2 => n695, ZN => n6243);
   U2472 : OAI222_X1 port map( A1 => n1007, A2 => n635, B1 => n1039, B2 => n632
                           , C1 => n975, C2 => n629, ZN => n6274);
   U2473 : OAI222_X1 port map( A1 => n303, A2 => n1413, B1 => n335, B2 => n1410
                           , C1 => n271, C2 => n1407, ZN => n4800);
   U2474 : OAI222_X1 port map( A1 => n1007, A2 => n1347, B1 => n1039, B2 => 
                           n1344, C1 => n975, C2 => n1341, ZN => n4831);
   U2475 : OAI222_X1 port map( A1 => n302, A2 => n701, B1 => n334, B2 => n698, 
                           C1 => n270, C2 => n695, ZN => n6202);
   U2476 : OAI222_X1 port map( A1 => n1006, A2 => n635, B1 => n1038, B2 => n632
                           , C1 => n974, C2 => n629, ZN => n6211);
   U2477 : OAI222_X1 port map( A1 => n302, A2 => n1413, B1 => n334, B2 => n1410
                           , C1 => n270, C2 => n1407, ZN => n4759);
   U2478 : OAI222_X1 port map( A1 => n1006, A2 => n1347, B1 => n1038, B2 => 
                           n1344, C1 => n974, C2 => n1341, ZN => n4768);
   U2479 : OAI222_X1 port map( A1 => n301, A2 => n701, B1 => n333, B2 => n698, 
                           C1 => n269, C2 => n695, ZN => n6161);
   U2480 : OAI222_X1 port map( A1 => n1005, A2 => n635, B1 => n1037, B2 => n632
                           , C1 => n973, C2 => n629, ZN => n6170);
   U2481 : OAI222_X1 port map( A1 => n301, A2 => n1413, B1 => n333, B2 => n1410
                           , C1 => n269, C2 => n1407, ZN => n4718);
   U2482 : OAI222_X1 port map( A1 => n1005, A2 => n1347, B1 => n1037, B2 => 
                           n1344, C1 => n973, C2 => n1341, ZN => n4727);
   U2483 : OAI222_X1 port map( A1 => n300, A2 => n701, B1 => n332, B2 => n698, 
                           C1 => n268, C2 => n695, ZN => n6120);
   U2484 : OAI222_X1 port map( A1 => n1004, A2 => n635, B1 => n1036, B2 => n632
                           , C1 => n972, C2 => n629, ZN => n6129);
   U2485 : OAI222_X1 port map( A1 => n300, A2 => n1413, B1 => n332, B2 => n1410
                           , C1 => n268, C2 => n1407, ZN => n4677);
   U2486 : OAI222_X1 port map( A1 => n1004, A2 => n1347, B1 => n1036, B2 => 
                           n1344, C1 => n972, C2 => n1341, ZN => n4686);
   U2487 : OAI222_X1 port map( A1 => n299, A2 => n701, B1 => n331, B2 => n698, 
                           C1 => n267, C2 => n695, ZN => n6079);
   U2488 : OAI222_X1 port map( A1 => n1003, A2 => n635, B1 => n1035, B2 => n632
                           , C1 => n971, C2 => n629, ZN => n6088);
   U2489 : OAI222_X1 port map( A1 => n299, A2 => n1413, B1 => n331, B2 => n1410
                           , C1 => n267, C2 => n1407, ZN => n4636);
   U2490 : OAI222_X1 port map( A1 => n1003, A2 => n1347, B1 => n1035, B2 => 
                           n1344, C1 => n971, C2 => n1341, ZN => n4645);
   U2491 : OAI222_X1 port map( A1 => n298, A2 => n701, B1 => n330, B2 => n698, 
                           C1 => n266, C2 => n695, ZN => n6038);
   U2492 : OAI222_X1 port map( A1 => n1002, A2 => n635, B1 => n1034, B2 => n632
                           , C1 => n970, C2 => n629, ZN => n6047);
   U2493 : OAI222_X1 port map( A1 => n298, A2 => n1413, B1 => n330, B2 => n1410
                           , C1 => n266, C2 => n1407, ZN => n4595);
   U2494 : OAI222_X1 port map( A1 => n1002, A2 => n1347, B1 => n1034, B2 => 
                           n1344, C1 => n970, C2 => n1341, ZN => n4604);
   U2495 : OAI222_X1 port map( A1 => n297, A2 => n701, B1 => n329, B2 => n698, 
                           C1 => n265, C2 => n695, ZN => n5997);
   U2496 : OAI222_X1 port map( A1 => n1001, A2 => n635, B1 => n1033, B2 => n632
                           , C1 => n969, C2 => n629, ZN => n6006);
   U2497 : OAI222_X1 port map( A1 => n297, A2 => n1413, B1 => n329, B2 => n1410
                           , C1 => n265, C2 => n1407, ZN => n4554);
   U2498 : OAI222_X1 port map( A1 => n1001, A2 => n1347, B1 => n1033, B2 => 
                           n1344, C1 => n969, C2 => n1341, ZN => n4563);
   U2499 : OAI222_X1 port map( A1 => n296, A2 => n701, B1 => n328, B2 => n698, 
                           C1 => n264, C2 => n695, ZN => n5956);
   U2500 : OAI222_X1 port map( A1 => n1000, A2 => n635, B1 => n1032, B2 => n632
                           , C1 => n968, C2 => n629, ZN => n5965);
   U2501 : OAI222_X1 port map( A1 => n296, A2 => n1413, B1 => n328, B2 => n1410
                           , C1 => n264, C2 => n1407, ZN => n4513);
   U2502 : OAI222_X1 port map( A1 => n1000, A2 => n1347, B1 => n1032, B2 => 
                           n1344, C1 => n968, C2 => n1341, ZN => n4522);
   U2503 : OAI222_X1 port map( A1 => n295, A2 => n701, B1 => n327, B2 => n698, 
                           C1 => n263, C2 => n695, ZN => n5915);
   U2504 : OAI222_X1 port map( A1 => n999, A2 => n635, B1 => n1031, B2 => n632,
                           C1 => n967, C2 => n629, ZN => n5924);
   U2505 : OAI222_X1 port map( A1 => n295, A2 => n1413, B1 => n327, B2 => n1410
                           , C1 => n263, C2 => n1407, ZN => n4472);
   U2506 : OAI222_X1 port map( A1 => n999, A2 => n1347, B1 => n1031, B2 => 
                           n1344, C1 => n967, C2 => n1341, ZN => n4481);
   U2507 : OAI222_X1 port map( A1 => n294, A2 => n701, B1 => n326, B2 => n698, 
                           C1 => n262, C2 => n695, ZN => n5874);
   U2508 : OAI222_X1 port map( A1 => n998, A2 => n635, B1 => n1030, B2 => n632,
                           C1 => n966, C2 => n629, ZN => n5883);
   U2509 : OAI222_X1 port map( A1 => n294, A2 => n1413, B1 => n326, B2 => n1410
                           , C1 => n262, C2 => n1407, ZN => n4431);
   U2510 : OAI222_X1 port map( A1 => n998, A2 => n1347, B1 => n1030, B2 => 
                           n1344, C1 => n966, C2 => n1341, ZN => n4440);
   U2511 : OAI222_X1 port map( A1 => n293, A2 => n701, B1 => n325, B2 => n698, 
                           C1 => n261, C2 => n695, ZN => n5833);
   U2512 : OAI222_X1 port map( A1 => n997, A2 => n635, B1 => n1029, B2 => n632,
                           C1 => n965, C2 => n629, ZN => n5842);
   U2513 : OAI222_X1 port map( A1 => n293, A2 => n1413, B1 => n325, B2 => n1410
                           , C1 => n261, C2 => n1407, ZN => n4390);
   U2514 : OAI222_X1 port map( A1 => n997, A2 => n1347, B1 => n1029, B2 => 
                           n1344, C1 => n965, C2 => n1341, ZN => n4399);
   U2515 : OAI222_X1 port map( A1 => n292, A2 => n701, B1 => n324, B2 => n698, 
                           C1 => n260, C2 => n695, ZN => n5792);
   U2516 : OAI222_X1 port map( A1 => n996, A2 => n635, B1 => n1028, B2 => n632,
                           C1 => n964, C2 => n629, ZN => n5801);
   U2517 : OAI222_X1 port map( A1 => n292, A2 => n1413, B1 => n324, B2 => n1410
                           , C1 => n260, C2 => n1407, ZN => n4349);
   U2518 : OAI222_X1 port map( A1 => n996, A2 => n1347, B1 => n1028, B2 => 
                           n1344, C1 => n964, C2 => n1341, ZN => n4358);
   U2519 : OAI222_X1 port map( A1 => n291, A2 => n702, B1 => n323, B2 => n699, 
                           C1 => n259, C2 => n696, ZN => n5751);
   U2520 : OAI222_X1 port map( A1 => n995, A2 => n636, B1 => n1027, B2 => n633,
                           C1 => n963, C2 => n630, ZN => n5760);
   U2521 : OAI222_X1 port map( A1 => n291, A2 => n1414, B1 => n323, B2 => n1411
                           , C1 => n259, C2 => n1408, ZN => n4308);
   U2522 : OAI222_X1 port map( A1 => n995, A2 => n1348, B1 => n1027, B2 => 
                           n1345, C1 => n963, C2 => n1342, ZN => n4317);
   U2523 : OAI222_X1 port map( A1 => n290, A2 => n702, B1 => n322, B2 => n699, 
                           C1 => n258, C2 => n696, ZN => n5710);
   U2524 : OAI222_X1 port map( A1 => n994, A2 => n636, B1 => n1026, B2 => n633,
                           C1 => n962, C2 => n630, ZN => n5719);
   U2525 : OAI222_X1 port map( A1 => n290, A2 => n1414, B1 => n322, B2 => n1411
                           , C1 => n258, C2 => n1408, ZN => n4267);
   U2526 : OAI222_X1 port map( A1 => n994, A2 => n1348, B1 => n1026, B2 => 
                           n1345, C1 => n962, C2 => n1342, ZN => n4276);
   U2527 : OAI222_X1 port map( A1 => n289, A2 => n702, B1 => n321, B2 => n699, 
                           C1 => n257, C2 => n696, ZN => n5669);
   U2528 : OAI222_X1 port map( A1 => n993, A2 => n636, B1 => n1025, B2 => n633,
                           C1 => n961, C2 => n630, ZN => n5678);
   U2529 : OAI222_X1 port map( A1 => n289, A2 => n1414, B1 => n321, B2 => n1411
                           , C1 => n257, C2 => n1408, ZN => n4226);
   U2530 : OAI222_X1 port map( A1 => n993, A2 => n1348, B1 => n1025, B2 => 
                           n1345, C1 => n961, C2 => n1342, ZN => n4235);
   U2531 : OAI222_X1 port map( A1 => n288, A2 => n702, B1 => n320, B2 => n699, 
                           C1 => n256, C2 => n696, ZN => n5628);
   U2532 : OAI222_X1 port map( A1 => n992, A2 => n636, B1 => n1024, B2 => n633,
                           C1 => n960, C2 => n630, ZN => n5637);
   U2533 : OAI222_X1 port map( A1 => n288, A2 => n1414, B1 => n320, B2 => n1411
                           , C1 => n256, C2 => n1408, ZN => n4185);
   U2534 : OAI222_X1 port map( A1 => n992, A2 => n1348, B1 => n1024, B2 => 
                           n1345, C1 => n960, C2 => n1342, ZN => n4194);
   U2535 : OAI222_X1 port map( A1 => n287, A2 => n702, B1 => n319, B2 => n699, 
                           C1 => n255, C2 => n696, ZN => n5587);
   U2536 : OAI222_X1 port map( A1 => n991, A2 => n636, B1 => n1023, B2 => n633,
                           C1 => n959, C2 => n630, ZN => n5596);
   U2537 : OAI222_X1 port map( A1 => n287, A2 => n1414, B1 => n319, B2 => n1411
                           , C1 => n255, C2 => n1408, ZN => n4144);
   U2538 : OAI222_X1 port map( A1 => n991, A2 => n1348, B1 => n1023, B2 => 
                           n1345, C1 => n959, C2 => n1342, ZN => n4153);
   U2539 : OAI222_X1 port map( A1 => n286, A2 => n702, B1 => n318, B2 => n699, 
                           C1 => n254, C2 => n696, ZN => n5546);
   U2540 : OAI222_X1 port map( A1 => n990, A2 => n636, B1 => n1022, B2 => n633,
                           C1 => n958, C2 => n630, ZN => n5555);
   U2541 : OAI222_X1 port map( A1 => n286, A2 => n1414, B1 => n318, B2 => n1411
                           , C1 => n254, C2 => n1408, ZN => n4103);
   U2542 : OAI222_X1 port map( A1 => n990, A2 => n1348, B1 => n1022, B2 => 
                           n1345, C1 => n958, C2 => n1342, ZN => n4112);
   U2543 : OAI222_X1 port map( A1 => n285, A2 => n702, B1 => n317, B2 => n699, 
                           C1 => n253, C2 => n696, ZN => n5505);
   U2544 : OAI222_X1 port map( A1 => n989, A2 => n636, B1 => n1021, B2 => n633,
                           C1 => n957, C2 => n630, ZN => n5514);
   U2545 : OAI222_X1 port map( A1 => n285, A2 => n1414, B1 => n317, B2 => n1411
                           , C1 => n253, C2 => n1408, ZN => n4062);
   U2546 : OAI222_X1 port map( A1 => n989, A2 => n1348, B1 => n1021, B2 => 
                           n1345, C1 => n957, C2 => n1342, ZN => n4071);
   U2547 : OAI222_X1 port map( A1 => n284, A2 => n702, B1 => n316, B2 => n699, 
                           C1 => n252, C2 => n696, ZN => n5464);
   U2548 : OAI222_X1 port map( A1 => n988, A2 => n636, B1 => n1020, B2 => n633,
                           C1 => n956, C2 => n630, ZN => n5473);
   U2549 : OAI222_X1 port map( A1 => n284, A2 => n1414, B1 => n316, B2 => n1411
                           , C1 => n252, C2 => n1408, ZN => n4021);
   U2550 : OAI222_X1 port map( A1 => n988, A2 => n1348, B1 => n1020, B2 => 
                           n1345, C1 => n956, C2 => n1342, ZN => n4030);
   U2551 : OAI222_X1 port map( A1 => n283, A2 => n702, B1 => n315, B2 => n699, 
                           C1 => n251, C2 => n696, ZN => n5423);
   U2552 : OAI222_X1 port map( A1 => n987, A2 => n636, B1 => n1019, B2 => n633,
                           C1 => n955, C2 => n630, ZN => n5432);
   U2553 : OAI222_X1 port map( A1 => n283, A2 => n1414, B1 => n315, B2 => n1411
                           , C1 => n251, C2 => n1408, ZN => n3980);
   U2554 : OAI222_X1 port map( A1 => n987, A2 => n1348, B1 => n1019, B2 => 
                           n1345, C1 => n955, C2 => n1342, ZN => n3989);
   U2555 : OAI222_X1 port map( A1 => n282, A2 => n702, B1 => n314, B2 => n699, 
                           C1 => n250, C2 => n696, ZN => n5382);
   U2556 : OAI222_X1 port map( A1 => n986, A2 => n636, B1 => n1018, B2 => n633,
                           C1 => n954, C2 => n630, ZN => n5391);
   U2557 : OAI222_X1 port map( A1 => n282, A2 => n1414, B1 => n314, B2 => n1411
                           , C1 => n250, C2 => n1408, ZN => n3939);
   U2558 : OAI222_X1 port map( A1 => n986, A2 => n1348, B1 => n1018, B2 => 
                           n1345, C1 => n954, C2 => n1342, ZN => n3948);
   U2559 : OAI222_X1 port map( A1 => n281, A2 => n702, B1 => n313, B2 => n699, 
                           C1 => n249, C2 => n696, ZN => n5341);
   U2560 : OAI222_X1 port map( A1 => n985, A2 => n636, B1 => n1017, B2 => n633,
                           C1 => n953, C2 => n630, ZN => n5350);
   U2561 : OAI222_X1 port map( A1 => n281, A2 => n1414, B1 => n313, B2 => n1411
                           , C1 => n249, C2 => n1408, ZN => n3898);
   U2562 : OAI222_X1 port map( A1 => n985, A2 => n1348, B1 => n1017, B2 => 
                           n1345, C1 => n953, C2 => n1342, ZN => n3907);
   U2563 : OAI222_X1 port map( A1 => n280, A2 => n702, B1 => n312, B2 => n699, 
                           C1 => n248, C2 => n696, ZN => n5300);
   U2564 : OAI222_X1 port map( A1 => n984, A2 => n636, B1 => n1016, B2 => n633,
                           C1 => n952, C2 => n630, ZN => n5309);
   U2565 : OAI222_X1 port map( A1 => n280, A2 => n1414, B1 => n312, B2 => n1411
                           , C1 => n248, C2 => n1408, ZN => n3857);
   U2566 : OAI222_X1 port map( A1 => n984, A2 => n1348, B1 => n1016, B2 => 
                           n1345, C1 => n952, C2 => n1342, ZN => n3866);
   U2567 : OAI222_X1 port map( A1 => n279, A2 => n703, B1 => n311, B2 => n700, 
                           C1 => n247, C2 => n697, ZN => n5259);
   U2568 : OAI222_X1 port map( A1 => n983, A2 => n637, B1 => n1015, B2 => n634,
                           C1 => n951, C2 => n631, ZN => n5268);
   U2569 : OAI222_X1 port map( A1 => n279, A2 => n1415, B1 => n311, B2 => n1412
                           , C1 => n247, C2 => n1409, ZN => n3816);
   U2570 : OAI222_X1 port map( A1 => n983, A2 => n1349, B1 => n1015, B2 => 
                           n1346, C1 => n951, C2 => n1343, ZN => n3825);
   U2571 : OAI222_X1 port map( A1 => n278, A2 => n703, B1 => n310, B2 => n700, 
                           C1 => n246, C2 => n697, ZN => n5218);
   U2572 : OAI222_X1 port map( A1 => n982, A2 => n637, B1 => n1014, B2 => n634,
                           C1 => n950, C2 => n631, ZN => n5227);
   U2573 : OAI222_X1 port map( A1 => n278, A2 => n1415, B1 => n310, B2 => n1412
                           , C1 => n246, C2 => n1409, ZN => n3775);
   U2574 : OAI222_X1 port map( A1 => n982, A2 => n1349, B1 => n1014, B2 => 
                           n1346, C1 => n950, C2 => n1343, ZN => n3784);
   U2575 : OAI222_X1 port map( A1 => n277, A2 => n703, B1 => n309, B2 => n700, 
                           C1 => n245, C2 => n697, ZN => n5177);
   U2576 : OAI222_X1 port map( A1 => n981, A2 => n637, B1 => n1013, B2 => n634,
                           C1 => n949, C2 => n631, ZN => n5186);
   U2577 : OAI222_X1 port map( A1 => n277, A2 => n1415, B1 => n309, B2 => n1412
                           , C1 => n245, C2 => n1409, ZN => n3734);
   U2578 : OAI222_X1 port map( A1 => n981, A2 => n1349, B1 => n1013, B2 => 
                           n1346, C1 => n949, C2 => n1343, ZN => n3743);
   U2579 : OAI222_X1 port map( A1 => n276, A2 => n703, B1 => n308, B2 => n700, 
                           C1 => n244, C2 => n697, ZN => n5136);
   U2580 : OAI222_X1 port map( A1 => n980, A2 => n637, B1 => n1012, B2 => n634,
                           C1 => n948, C2 => n631, ZN => n5145);
   U2581 : OAI222_X1 port map( A1 => n276, A2 => n1415, B1 => n308, B2 => n1412
                           , C1 => n244, C2 => n1409, ZN => n3693);
   U2582 : OAI222_X1 port map( A1 => n980, A2 => n1349, B1 => n1012, B2 => 
                           n1346, C1 => n948, C2 => n1343, ZN => n3702);
   U2583 : OAI222_X1 port map( A1 => n275, A2 => n703, B1 => n307, B2 => n700, 
                           C1 => n243, C2 => n697, ZN => n5095);
   U2584 : OAI222_X1 port map( A1 => n979, A2 => n637, B1 => n1011, B2 => n634,
                           C1 => n947, C2 => n631, ZN => n5104);
   U2585 : OAI222_X1 port map( A1 => n275, A2 => n1415, B1 => n307, B2 => n1412
                           , C1 => n243, C2 => n1409, ZN => n3652);
   U2586 : OAI222_X1 port map( A1 => n979, A2 => n1349, B1 => n1011, B2 => 
                           n1346, C1 => n947, C2 => n1343, ZN => n3661);
   U2587 : OAI222_X1 port map( A1 => n274, A2 => n703, B1 => n306, B2 => n700, 
                           C1 => n242, C2 => n697, ZN => n5054);
   U2588 : OAI222_X1 port map( A1 => n978, A2 => n637, B1 => n1010, B2 => n634,
                           C1 => n946, C2 => n631, ZN => n5063);
   U2589 : OAI222_X1 port map( A1 => n274, A2 => n1415, B1 => n306, B2 => n1412
                           , C1 => n242, C2 => n1409, ZN => n3611);
   U2590 : OAI222_X1 port map( A1 => n978, A2 => n1349, B1 => n1010, B2 => 
                           n1346, C1 => n946, C2 => n1343, ZN => n3620);
   U2591 : OAI222_X1 port map( A1 => n273, A2 => n703, B1 => n305, B2 => n700, 
                           C1 => n241, C2 => n697, ZN => n5013);
   U2592 : OAI222_X1 port map( A1 => n977, A2 => n637, B1 => n1009, B2 => n634,
                           C1 => n945, C2 => n631, ZN => n5022);
   U2593 : OAI222_X1 port map( A1 => n273, A2 => n1415, B1 => n305, B2 => n1412
                           , C1 => n241, C2 => n1409, ZN => n3570);
   U2594 : OAI222_X1 port map( A1 => n977, A2 => n1349, B1 => n1009, B2 => 
                           n1346, C1 => n945, C2 => n1343, ZN => n3579);
   U2595 : OAI222_X1 port map( A1 => n272, A2 => n703, B1 => n304, B2 => n700, 
                           C1 => n240, C2 => n697, ZN => n4884);
   U2596 : OAI222_X1 port map( A1 => n976, A2 => n637, B1 => n1008, B2 => n634,
                           C1 => n944, C2 => n631, ZN => n4915);
   U2597 : OAI222_X1 port map( A1 => n272, A2 => n1415, B1 => n304, B2 => n1412
                           , C1 => n240, C2 => n1409, ZN => n3441);
   U2598 : OAI222_X1 port map( A1 => n976, A2 => n1349, B1 => n1008, B2 => 
                           n1346, C1 => n944, C2 => n1343, ZN => n3472);
   U2599 : OAI222_X1 port map( A1 => n399, A2 => n692, B1 => n431, B2 => n689, 
                           C1 => n367, C2 => n686, ZN => n6242);
   U2600 : OAI222_X1 port map( A1 => n1103, A2 => n626, B1 => n1135, B2 => n623
                           , C1 => n1071, C2 => n620, ZN => n6273);
   U2601 : OAI222_X1 port map( A1 => n399, A2 => n1404, B1 => n431, B2 => n1401
                           , C1 => n367, C2 => n1398, ZN => n4799);
   U2602 : OAI222_X1 port map( A1 => n1103, A2 => n1338, B1 => n1135, B2 => 
                           n1335, C1 => n1071, C2 => n1332, ZN => n4830);
   U2603 : OAI222_X1 port map( A1 => n398, A2 => n692, B1 => n430, B2 => n689, 
                           C1 => n366, C2 => n686, ZN => n6201);
   U2604 : OAI222_X1 port map( A1 => n1102, A2 => n626, B1 => n1134, B2 => n623
                           , C1 => n1070, C2 => n620, ZN => n6210);
   U2605 : OAI222_X1 port map( A1 => n398, A2 => n1404, B1 => n430, B2 => n1401
                           , C1 => n366, C2 => n1398, ZN => n4758);
   U2606 : OAI222_X1 port map( A1 => n1102, A2 => n1338, B1 => n1134, B2 => 
                           n1335, C1 => n1070, C2 => n1332, ZN => n4767);
   U2607 : OAI222_X1 port map( A1 => n397, A2 => n692, B1 => n429, B2 => n689, 
                           C1 => n365, C2 => n686, ZN => n6160);
   U2608 : OAI222_X1 port map( A1 => n1101, A2 => n626, B1 => n1133, B2 => n623
                           , C1 => n1069, C2 => n620, ZN => n6169);
   U2609 : OAI222_X1 port map( A1 => n397, A2 => n1404, B1 => n429, B2 => n1401
                           , C1 => n365, C2 => n1398, ZN => n4717);
   U2610 : OAI222_X1 port map( A1 => n1101, A2 => n1338, B1 => n1133, B2 => 
                           n1335, C1 => n1069, C2 => n1332, ZN => n4726);
   U2611 : OAI222_X1 port map( A1 => n396, A2 => n692, B1 => n428, B2 => n689, 
                           C1 => n364, C2 => n686, ZN => n6119);
   U2612 : OAI222_X1 port map( A1 => n1100, A2 => n626, B1 => n1132, B2 => n623
                           , C1 => n1068, C2 => n620, ZN => n6128);
   U2613 : OAI222_X1 port map( A1 => n396, A2 => n1404, B1 => n428, B2 => n1401
                           , C1 => n364, C2 => n1398, ZN => n4676);
   U2614 : OAI222_X1 port map( A1 => n1100, A2 => n1338, B1 => n1132, B2 => 
                           n1335, C1 => n1068, C2 => n1332, ZN => n4685);
   U2615 : OAI222_X1 port map( A1 => n395, A2 => n692, B1 => n427, B2 => n689, 
                           C1 => n363, C2 => n686, ZN => n6078);
   U2616 : OAI222_X1 port map( A1 => n1099, A2 => n626, B1 => n1131, B2 => n623
                           , C1 => n1067, C2 => n620, ZN => n6087);
   U2617 : OAI222_X1 port map( A1 => n395, A2 => n1404, B1 => n427, B2 => n1401
                           , C1 => n363, C2 => n1398, ZN => n4635);
   U2618 : OAI222_X1 port map( A1 => n1099, A2 => n1338, B1 => n1131, B2 => 
                           n1335, C1 => n1067, C2 => n1332, ZN => n4644);
   U2619 : OAI222_X1 port map( A1 => n394, A2 => n692, B1 => n426, B2 => n689, 
                           C1 => n362, C2 => n686, ZN => n6037);
   U2620 : OAI222_X1 port map( A1 => n1098, A2 => n626, B1 => n1130, B2 => n623
                           , C1 => n1066, C2 => n620, ZN => n6046);
   U2621 : OAI222_X1 port map( A1 => n394, A2 => n1404, B1 => n426, B2 => n1401
                           , C1 => n362, C2 => n1398, ZN => n4594);
   U2622 : OAI222_X1 port map( A1 => n1098, A2 => n1338, B1 => n1130, B2 => 
                           n1335, C1 => n1066, C2 => n1332, ZN => n4603);
   U2623 : OAI222_X1 port map( A1 => n393, A2 => n692, B1 => n425, B2 => n689, 
                           C1 => n361, C2 => n686, ZN => n5996);
   U2624 : OAI222_X1 port map( A1 => n1097, A2 => n626, B1 => n1129, B2 => n623
                           , C1 => n1065, C2 => n620, ZN => n6005);
   U2625 : OAI222_X1 port map( A1 => n393, A2 => n1404, B1 => n425, B2 => n1401
                           , C1 => n361, C2 => n1398, ZN => n4553);
   U2626 : OAI222_X1 port map( A1 => n1097, A2 => n1338, B1 => n1129, B2 => 
                           n1335, C1 => n1065, C2 => n1332, ZN => n4562);
   U2627 : OAI222_X1 port map( A1 => n392, A2 => n692, B1 => n424, B2 => n689, 
                           C1 => n360, C2 => n686, ZN => n5955);
   U2628 : OAI222_X1 port map( A1 => n1096, A2 => n626, B1 => n1128, B2 => n623
                           , C1 => n1064, C2 => n620, ZN => n5964);
   U2629 : OAI222_X1 port map( A1 => n392, A2 => n1404, B1 => n424, B2 => n1401
                           , C1 => n360, C2 => n1398, ZN => n4512);
   U2630 : OAI222_X1 port map( A1 => n1096, A2 => n1338, B1 => n1128, B2 => 
                           n1335, C1 => n1064, C2 => n1332, ZN => n4521);
   U2631 : OAI222_X1 port map( A1 => n391, A2 => n692, B1 => n423, B2 => n689, 
                           C1 => n359, C2 => n686, ZN => n5914);
   U2632 : OAI222_X1 port map( A1 => n1095, A2 => n626, B1 => n1127, B2 => n623
                           , C1 => n1063, C2 => n620, ZN => n5923);
   U2633 : OAI222_X1 port map( A1 => n391, A2 => n1404, B1 => n423, B2 => n1401
                           , C1 => n359, C2 => n1398, ZN => n4471);
   U2634 : OAI222_X1 port map( A1 => n1095, A2 => n1338, B1 => n1127, B2 => 
                           n1335, C1 => n1063, C2 => n1332, ZN => n4480);
   U2635 : OAI222_X1 port map( A1 => n390, A2 => n692, B1 => n422, B2 => n689, 
                           C1 => n358, C2 => n686, ZN => n5873);
   U2636 : OAI222_X1 port map( A1 => n1094, A2 => n626, B1 => n1126, B2 => n623
                           , C1 => n1062, C2 => n620, ZN => n5882);
   U2637 : OAI222_X1 port map( A1 => n390, A2 => n1404, B1 => n422, B2 => n1401
                           , C1 => n358, C2 => n1398, ZN => n4430);
   U2638 : OAI222_X1 port map( A1 => n1094, A2 => n1338, B1 => n1126, B2 => 
                           n1335, C1 => n1062, C2 => n1332, ZN => n4439);
   U2639 : OAI222_X1 port map( A1 => n389, A2 => n692, B1 => n421, B2 => n689, 
                           C1 => n357, C2 => n686, ZN => n5832);
   U2640 : OAI222_X1 port map( A1 => n1093, A2 => n626, B1 => n1125, B2 => n623
                           , C1 => n1061, C2 => n620, ZN => n5841);
   U2641 : OAI222_X1 port map( A1 => n389, A2 => n1404, B1 => n421, B2 => n1401
                           , C1 => n357, C2 => n1398, ZN => n4389);
   U2642 : OAI222_X1 port map( A1 => n1093, A2 => n1338, B1 => n1125, B2 => 
                           n1335, C1 => n1061, C2 => n1332, ZN => n4398);
   U2643 : OAI222_X1 port map( A1 => n388, A2 => n692, B1 => n420, B2 => n689, 
                           C1 => n356, C2 => n686, ZN => n5791);
   U2644 : OAI222_X1 port map( A1 => n1092, A2 => n626, B1 => n1124, B2 => n623
                           , C1 => n1060, C2 => n620, ZN => n5800);
   U2645 : OAI222_X1 port map( A1 => n388, A2 => n1404, B1 => n420, B2 => n1401
                           , C1 => n356, C2 => n1398, ZN => n4348);
   U2646 : OAI222_X1 port map( A1 => n1092, A2 => n1338, B1 => n1124, B2 => 
                           n1335, C1 => n1060, C2 => n1332, ZN => n4357);
   U2647 : OAI222_X1 port map( A1 => n387, A2 => n693, B1 => n419, B2 => n690, 
                           C1 => n355, C2 => n687, ZN => n5750);
   U2648 : OAI222_X1 port map( A1 => n1091, A2 => n627, B1 => n1123, B2 => n624
                           , C1 => n1059, C2 => n621, ZN => n5759);
   U2649 : OAI222_X1 port map( A1 => n387, A2 => n1405, B1 => n419, B2 => n1402
                           , C1 => n355, C2 => n1399, ZN => n4307);
   U2650 : OAI222_X1 port map( A1 => n1091, A2 => n1339, B1 => n1123, B2 => 
                           n1336, C1 => n1059, C2 => n1333, ZN => n4316);
   U2651 : OAI222_X1 port map( A1 => n386, A2 => n693, B1 => n418, B2 => n690, 
                           C1 => n354, C2 => n687, ZN => n5709);
   U2652 : OAI222_X1 port map( A1 => n1090, A2 => n627, B1 => n1122, B2 => n624
                           , C1 => n1058, C2 => n621, ZN => n5718);
   U2653 : OAI222_X1 port map( A1 => n386, A2 => n1405, B1 => n418, B2 => n1402
                           , C1 => n354, C2 => n1399, ZN => n4266);
   U2654 : OAI222_X1 port map( A1 => n1090, A2 => n1339, B1 => n1122, B2 => 
                           n1336, C1 => n1058, C2 => n1333, ZN => n4275);
   U2655 : OAI222_X1 port map( A1 => n385, A2 => n693, B1 => n417, B2 => n690, 
                           C1 => n353, C2 => n687, ZN => n5668);
   U2656 : OAI222_X1 port map( A1 => n1089, A2 => n627, B1 => n1121, B2 => n624
                           , C1 => n1057, C2 => n621, ZN => n5677);
   U2657 : OAI222_X1 port map( A1 => n385, A2 => n1405, B1 => n417, B2 => n1402
                           , C1 => n353, C2 => n1399, ZN => n4225);
   U2658 : OAI222_X1 port map( A1 => n1089, A2 => n1339, B1 => n1121, B2 => 
                           n1336, C1 => n1057, C2 => n1333, ZN => n4234);
   U2659 : OAI222_X1 port map( A1 => n384, A2 => n693, B1 => n416, B2 => n690, 
                           C1 => n352, C2 => n687, ZN => n5627);
   U2660 : OAI222_X1 port map( A1 => n1088, A2 => n627, B1 => n1120, B2 => n624
                           , C1 => n1056, C2 => n621, ZN => n5636);
   U2661 : OAI222_X1 port map( A1 => n384, A2 => n1405, B1 => n416, B2 => n1402
                           , C1 => n352, C2 => n1399, ZN => n4184);
   U2662 : OAI222_X1 port map( A1 => n1088, A2 => n1339, B1 => n1120, B2 => 
                           n1336, C1 => n1056, C2 => n1333, ZN => n4193);
   U2663 : OAI222_X1 port map( A1 => n383, A2 => n693, B1 => n415, B2 => n690, 
                           C1 => n351, C2 => n687, ZN => n5586);
   U2664 : OAI222_X1 port map( A1 => n1087, A2 => n627, B1 => n1119, B2 => n624
                           , C1 => n1055, C2 => n621, ZN => n5595);
   U2665 : OAI222_X1 port map( A1 => n383, A2 => n1405, B1 => n415, B2 => n1402
                           , C1 => n351, C2 => n1399, ZN => n4143);
   U2666 : OAI222_X1 port map( A1 => n1087, A2 => n1339, B1 => n1119, B2 => 
                           n1336, C1 => n1055, C2 => n1333, ZN => n4152);
   U2667 : OAI222_X1 port map( A1 => n382, A2 => n693, B1 => n414, B2 => n690, 
                           C1 => n350, C2 => n687, ZN => n5545);
   U2668 : OAI222_X1 port map( A1 => n1086, A2 => n627, B1 => n1118, B2 => n624
                           , C1 => n1054, C2 => n621, ZN => n5554);
   U2669 : OAI222_X1 port map( A1 => n382, A2 => n1405, B1 => n414, B2 => n1402
                           , C1 => n350, C2 => n1399, ZN => n4102);
   U2670 : OAI222_X1 port map( A1 => n1086, A2 => n1339, B1 => n1118, B2 => 
                           n1336, C1 => n1054, C2 => n1333, ZN => n4111);
   U2671 : OAI222_X1 port map( A1 => n381, A2 => n693, B1 => n413, B2 => n690, 
                           C1 => n349, C2 => n687, ZN => n5504);
   U2672 : OAI222_X1 port map( A1 => n1085, A2 => n627, B1 => n1117, B2 => n624
                           , C1 => n1053, C2 => n621, ZN => n5513);
   U2673 : OAI222_X1 port map( A1 => n381, A2 => n1405, B1 => n413, B2 => n1402
                           , C1 => n349, C2 => n1399, ZN => n4061);
   U2674 : OAI222_X1 port map( A1 => n1085, A2 => n1339, B1 => n1117, B2 => 
                           n1336, C1 => n1053, C2 => n1333, ZN => n4070);
   U2675 : OAI222_X1 port map( A1 => n380, A2 => n693, B1 => n412, B2 => n690, 
                           C1 => n348, C2 => n687, ZN => n5463);
   U2676 : OAI222_X1 port map( A1 => n1084, A2 => n627, B1 => n1116, B2 => n624
                           , C1 => n1052, C2 => n621, ZN => n5472);
   U2677 : OAI222_X1 port map( A1 => n380, A2 => n1405, B1 => n412, B2 => n1402
                           , C1 => n348, C2 => n1399, ZN => n4020);
   U2678 : OAI222_X1 port map( A1 => n1084, A2 => n1339, B1 => n1116, B2 => 
                           n1336, C1 => n1052, C2 => n1333, ZN => n4029);
   U2679 : OAI222_X1 port map( A1 => n379, A2 => n693, B1 => n411, B2 => n690, 
                           C1 => n347, C2 => n687, ZN => n5422);
   U2680 : OAI222_X1 port map( A1 => n1083, A2 => n627, B1 => n1115, B2 => n624
                           , C1 => n1051, C2 => n621, ZN => n5431);
   U2681 : OAI222_X1 port map( A1 => n379, A2 => n1405, B1 => n411, B2 => n1402
                           , C1 => n347, C2 => n1399, ZN => n3979);
   U2682 : OAI222_X1 port map( A1 => n1083, A2 => n1339, B1 => n1115, B2 => 
                           n1336, C1 => n1051, C2 => n1333, ZN => n3988);
   U2683 : OAI222_X1 port map( A1 => n378, A2 => n693, B1 => n410, B2 => n690, 
                           C1 => n346, C2 => n687, ZN => n5381);
   U2684 : OAI222_X1 port map( A1 => n1082, A2 => n627, B1 => n1114, B2 => n624
                           , C1 => n1050, C2 => n621, ZN => n5390);
   U2685 : OAI222_X1 port map( A1 => n378, A2 => n1405, B1 => n410, B2 => n1402
                           , C1 => n346, C2 => n1399, ZN => n3938);
   U2686 : OAI222_X1 port map( A1 => n1082, A2 => n1339, B1 => n1114, B2 => 
                           n1336, C1 => n1050, C2 => n1333, ZN => n3947);
   U2687 : OAI222_X1 port map( A1 => n377, A2 => n693, B1 => n409, B2 => n690, 
                           C1 => n345, C2 => n687, ZN => n5340);
   U2688 : OAI222_X1 port map( A1 => n1081, A2 => n627, B1 => n1113, B2 => n624
                           , C1 => n1049, C2 => n621, ZN => n5349);
   U2689 : OAI222_X1 port map( A1 => n377, A2 => n1405, B1 => n409, B2 => n1402
                           , C1 => n345, C2 => n1399, ZN => n3897);
   U2690 : OAI222_X1 port map( A1 => n1081, A2 => n1339, B1 => n1113, B2 => 
                           n1336, C1 => n1049, C2 => n1333, ZN => n3906);
   U2691 : OAI222_X1 port map( A1 => n376, A2 => n693, B1 => n408, B2 => n690, 
                           C1 => n344, C2 => n687, ZN => n5299);
   U2692 : OAI222_X1 port map( A1 => n1080, A2 => n627, B1 => n1112, B2 => n624
                           , C1 => n1048, C2 => n621, ZN => n5308);
   U2693 : OAI222_X1 port map( A1 => n376, A2 => n1405, B1 => n408, B2 => n1402
                           , C1 => n344, C2 => n1399, ZN => n3856);
   U2694 : OAI222_X1 port map( A1 => n1080, A2 => n1339, B1 => n1112, B2 => 
                           n1336, C1 => n1048, C2 => n1333, ZN => n3865);
   U2695 : OAI222_X1 port map( A1 => n375, A2 => n694, B1 => n407, B2 => n691, 
                           C1 => n343, C2 => n688, ZN => n5258);
   U2696 : OAI222_X1 port map( A1 => n1079, A2 => n628, B1 => n1111, B2 => n625
                           , C1 => n1047, C2 => n622, ZN => n5267);
   U2697 : OAI222_X1 port map( A1 => n375, A2 => n1406, B1 => n407, B2 => n1403
                           , C1 => n343, C2 => n1400, ZN => n3815);
   U2698 : OAI222_X1 port map( A1 => n1079, A2 => n1340, B1 => n1111, B2 => 
                           n1337, C1 => n1047, C2 => n1334, ZN => n3824);
   U2699 : OAI222_X1 port map( A1 => n374, A2 => n694, B1 => n406, B2 => n691, 
                           C1 => n342, C2 => n688, ZN => n5217);
   U2700 : OAI222_X1 port map( A1 => n1078, A2 => n628, B1 => n1110, B2 => n625
                           , C1 => n1046, C2 => n622, ZN => n5226);
   U2701 : OAI222_X1 port map( A1 => n374, A2 => n1406, B1 => n406, B2 => n1403
                           , C1 => n342, C2 => n1400, ZN => n3774);
   U2702 : OAI222_X1 port map( A1 => n1078, A2 => n1340, B1 => n1110, B2 => 
                           n1337, C1 => n1046, C2 => n1334, ZN => n3783);
   U2703 : OAI222_X1 port map( A1 => n373, A2 => n694, B1 => n405, B2 => n691, 
                           C1 => n341, C2 => n688, ZN => n5176);
   U2704 : OAI222_X1 port map( A1 => n1077, A2 => n628, B1 => n1109, B2 => n625
                           , C1 => n1045, C2 => n622, ZN => n5185);
   U2705 : OAI222_X1 port map( A1 => n373, A2 => n1406, B1 => n405, B2 => n1403
                           , C1 => n341, C2 => n1400, ZN => n3733);
   U2706 : OAI222_X1 port map( A1 => n1077, A2 => n1340, B1 => n1109, B2 => 
                           n1337, C1 => n1045, C2 => n1334, ZN => n3742);
   U2707 : OAI222_X1 port map( A1 => n372, A2 => n694, B1 => n404, B2 => n691, 
                           C1 => n340, C2 => n688, ZN => n5135);
   U2708 : OAI222_X1 port map( A1 => n1076, A2 => n628, B1 => n1108, B2 => n625
                           , C1 => n1044, C2 => n622, ZN => n5144);
   U2709 : OAI222_X1 port map( A1 => n372, A2 => n1406, B1 => n404, B2 => n1403
                           , C1 => n340, C2 => n1400, ZN => n3692);
   U2710 : OAI222_X1 port map( A1 => n1076, A2 => n1340, B1 => n1108, B2 => 
                           n1337, C1 => n1044, C2 => n1334, ZN => n3701);
   U2711 : OAI222_X1 port map( A1 => n371, A2 => n694, B1 => n403, B2 => n691, 
                           C1 => n339, C2 => n688, ZN => n5094);
   U2712 : OAI222_X1 port map( A1 => n1075, A2 => n628, B1 => n1107, B2 => n625
                           , C1 => n1043, C2 => n622, ZN => n5103);
   U2713 : OAI222_X1 port map( A1 => n371, A2 => n1406, B1 => n403, B2 => n1403
                           , C1 => n339, C2 => n1400, ZN => n3651);
   U2714 : OAI222_X1 port map( A1 => n1075, A2 => n1340, B1 => n1107, B2 => 
                           n1337, C1 => n1043, C2 => n1334, ZN => n3660);
   U2715 : OAI222_X1 port map( A1 => n370, A2 => n694, B1 => n402, B2 => n691, 
                           C1 => n338, C2 => n688, ZN => n5053);
   U2716 : OAI222_X1 port map( A1 => n1074, A2 => n628, B1 => n1106, B2 => n625
                           , C1 => n1042, C2 => n622, ZN => n5062);
   U2717 : OAI222_X1 port map( A1 => n370, A2 => n1406, B1 => n402, B2 => n1403
                           , C1 => n338, C2 => n1400, ZN => n3610);
   U2718 : OAI222_X1 port map( A1 => n1074, A2 => n1340, B1 => n1106, B2 => 
                           n1337, C1 => n1042, C2 => n1334, ZN => n3619);
   U2719 : OAI222_X1 port map( A1 => n369, A2 => n694, B1 => n401, B2 => n691, 
                           C1 => n337, C2 => n688, ZN => n5012);
   U2720 : OAI222_X1 port map( A1 => n1073, A2 => n628, B1 => n1105, B2 => n625
                           , C1 => n1041, C2 => n622, ZN => n5021);
   U2721 : OAI222_X1 port map( A1 => n369, A2 => n1406, B1 => n401, B2 => n1403
                           , C1 => n337, C2 => n1400, ZN => n3569);
   U2722 : OAI222_X1 port map( A1 => n1073, A2 => n1340, B1 => n1105, B2 => 
                           n1337, C1 => n1041, C2 => n1334, ZN => n3578);
   U2723 : OAI222_X1 port map( A1 => n368, A2 => n694, B1 => n400, B2 => n691, 
                           C1 => n336, C2 => n688, ZN => n4883);
   U2724 : OAI222_X1 port map( A1 => n1072, A2 => n628, B1 => n1104, B2 => n625
                           , C1 => n1040, C2 => n622, ZN => n4914);
   U2725 : OAI222_X1 port map( A1 => n368, A2 => n1406, B1 => n400, B2 => n1403
                           , C1 => n336, C2 => n1400, ZN => n3440);
   U2726 : OAI222_X1 port map( A1 => n1072, A2 => n1340, B1 => n1104, B2 => 
                           n1337, C1 => n1040, C2 => n1334, ZN => n3471);
   U2727 : AOI222_X1 port map( A1 => n79, A2 => REGISTERS_49_0_port, B1 => n78,
                           B2 => REGISTERS_51_0_port, C1 => n75, C2 => 
                           REGISTERS_50_0_port, ZN => n6288);
   U2728 : AOI222_X1 port map( A1 => n12, A2 => REGISTERS_82_0_port, B1 => n10,
                           B2 => REGISTERS_84_0_port, C1 => n6, C2 => 
                           REGISTERS_83_0_port, ZN => n6301);
   U2729 : AOI222_X1 port map( A1 => n1143, A2 => REGISTERS_49_0_port, B1 => 
                           n1142, B2 => REGISTERS_51_0_port, C1 => n1139, C2 =>
                           REGISTERS_50_0_port, ZN => n4845);
   U2730 : AOI222_X1 port map( A1 => n725, A2 => REGISTERS_82_0_port, B1 => 
                           n724, B2 => REGISTERS_84_0_port, C1 => n721, C2 => 
                           REGISTERS_83_0_port, ZN => n4858);
   U2731 : AOI222_X1 port map( A1 => n79, A2 => REGISTERS_49_1_port, B1 => n78,
                           B2 => REGISTERS_51_1_port, C1 => n75, C2 => 
                           REGISTERS_50_1_port, ZN => n6215);
   U2732 : AOI222_X1 port map( A1 => n12, A2 => REGISTERS_82_1_port, B1 => n10,
                           B2 => REGISTERS_84_1_port, C1 => n6, C2 => 
                           REGISTERS_83_1_port, ZN => n6224);
   U2733 : AOI222_X1 port map( A1 => n1143, A2 => REGISTERS_49_1_port, B1 => 
                           n1142, B2 => REGISTERS_51_1_port, C1 => n1139, C2 =>
                           REGISTERS_50_1_port, ZN => n4772);
   U2734 : AOI222_X1 port map( A1 => n725, A2 => REGISTERS_82_1_port, B1 => 
                           n724, B2 => REGISTERS_84_1_port, C1 => n721, C2 => 
                           REGISTERS_83_1_port, ZN => n4781);
   U2735 : AOI222_X1 port map( A1 => n79, A2 => REGISTERS_49_2_port, B1 => n78,
                           B2 => REGISTERS_51_2_port, C1 => n75, C2 => 
                           REGISTERS_50_2_port, ZN => n6174);
   U2736 : AOI222_X1 port map( A1 => n12, A2 => REGISTERS_82_2_port, B1 => n10,
                           B2 => REGISTERS_84_2_port, C1 => n6, C2 => 
                           REGISTERS_83_2_port, ZN => n6183);
   U2737 : AOI222_X1 port map( A1 => n1143, A2 => REGISTERS_49_2_port, B1 => 
                           n1142, B2 => REGISTERS_51_2_port, C1 => n1139, C2 =>
                           REGISTERS_50_2_port, ZN => n4731);
   U2738 : AOI222_X1 port map( A1 => n725, A2 => REGISTERS_82_2_port, B1 => 
                           n724, B2 => REGISTERS_84_2_port, C1 => n721, C2 => 
                           REGISTERS_83_2_port, ZN => n4740);
   U2739 : AOI222_X1 port map( A1 => n79, A2 => REGISTERS_49_3_port, B1 => n78,
                           B2 => REGISTERS_51_3_port, C1 => n75, C2 => 
                           REGISTERS_50_3_port, ZN => n6133);
   U2740 : AOI222_X1 port map( A1 => n12, A2 => REGISTERS_82_3_port, B1 => n10,
                           B2 => REGISTERS_84_3_port, C1 => n6, C2 => 
                           REGISTERS_83_3_port, ZN => n6142);
   U2741 : AOI222_X1 port map( A1 => n1143, A2 => REGISTERS_49_3_port, B1 => 
                           n1142, B2 => REGISTERS_51_3_port, C1 => n1139, C2 =>
                           REGISTERS_50_3_port, ZN => n4690);
   U2742 : AOI222_X1 port map( A1 => n725, A2 => REGISTERS_82_3_port, B1 => 
                           n724, B2 => REGISTERS_84_3_port, C1 => n721, C2 => 
                           REGISTERS_83_3_port, ZN => n4699);
   U2743 : AOI222_X1 port map( A1 => n79, A2 => REGISTERS_49_4_port, B1 => n78,
                           B2 => REGISTERS_51_4_port, C1 => n75, C2 => 
                           REGISTERS_50_4_port, ZN => n6092);
   U2744 : AOI222_X1 port map( A1 => n12, A2 => REGISTERS_82_4_port, B1 => n10,
                           B2 => REGISTERS_84_4_port, C1 => n6, C2 => 
                           REGISTERS_83_4_port, ZN => n6101);
   U2745 : AOI222_X1 port map( A1 => n1143, A2 => REGISTERS_49_4_port, B1 => 
                           n1142, B2 => REGISTERS_51_4_port, C1 => n1139, C2 =>
                           REGISTERS_50_4_port, ZN => n4649);
   U2746 : AOI222_X1 port map( A1 => n725, A2 => REGISTERS_82_4_port, B1 => 
                           n724, B2 => REGISTERS_84_4_port, C1 => n721, C2 => 
                           REGISTERS_83_4_port, ZN => n4658);
   U2747 : AOI222_X1 port map( A1 => n79, A2 => REGISTERS_49_5_port, B1 => n78,
                           B2 => REGISTERS_51_5_port, C1 => n75, C2 => 
                           REGISTERS_50_5_port, ZN => n6051);
   U2748 : AOI222_X1 port map( A1 => n12, A2 => REGISTERS_82_5_port, B1 => n10,
                           B2 => REGISTERS_84_5_port, C1 => n6, C2 => 
                           REGISTERS_83_5_port, ZN => n6060);
   U2749 : AOI222_X1 port map( A1 => n1143, A2 => REGISTERS_49_5_port, B1 => 
                           n1142, B2 => REGISTERS_51_5_port, C1 => n1139, C2 =>
                           REGISTERS_50_5_port, ZN => n4608);
   U2750 : AOI222_X1 port map( A1 => n725, A2 => REGISTERS_82_5_port, B1 => 
                           n724, B2 => REGISTERS_84_5_port, C1 => n721, C2 => 
                           REGISTERS_83_5_port, ZN => n4617);
   U2751 : AOI222_X1 port map( A1 => n79, A2 => REGISTERS_49_6_port, B1 => n78,
                           B2 => REGISTERS_51_6_port, C1 => n75, C2 => 
                           REGISTERS_50_6_port, ZN => n6010);
   U2752 : AOI222_X1 port map( A1 => n12, A2 => REGISTERS_82_6_port, B1 => n10,
                           B2 => REGISTERS_84_6_port, C1 => n6, C2 => 
                           REGISTERS_83_6_port, ZN => n6019);
   U2753 : AOI222_X1 port map( A1 => n1143, A2 => REGISTERS_49_6_port, B1 => 
                           n1142, B2 => REGISTERS_51_6_port, C1 => n1139, C2 =>
                           REGISTERS_50_6_port, ZN => n4567);
   U2754 : AOI222_X1 port map( A1 => n725, A2 => REGISTERS_82_6_port, B1 => 
                           n724, B2 => REGISTERS_84_6_port, C1 => n721, C2 => 
                           REGISTERS_83_6_port, ZN => n4576);
   U2755 : AOI222_X1 port map( A1 => n79, A2 => REGISTERS_49_7_port, B1 => n78,
                           B2 => REGISTERS_51_7_port, C1 => n75, C2 => 
                           REGISTERS_50_7_port, ZN => n5969);
   U2756 : AOI222_X1 port map( A1 => n12, A2 => REGISTERS_82_7_port, B1 => n10,
                           B2 => REGISTERS_84_7_port, C1 => n6, C2 => 
                           REGISTERS_83_7_port, ZN => n5978);
   U2757 : AOI222_X1 port map( A1 => n1143, A2 => REGISTERS_49_7_port, B1 => 
                           n1142, B2 => REGISTERS_51_7_port, C1 => n1139, C2 =>
                           REGISTERS_50_7_port, ZN => n4526);
   U2758 : AOI222_X1 port map( A1 => n725, A2 => REGISTERS_82_7_port, B1 => 
                           n724, B2 => REGISTERS_84_7_port, C1 => n721, C2 => 
                           REGISTERS_83_7_port, ZN => n4535);
   U2759 : AOI222_X1 port map( A1 => n79, A2 => REGISTERS_49_8_port, B1 => n77,
                           B2 => REGISTERS_51_8_port, C1 => n74, C2 => 
                           REGISTERS_50_8_port, ZN => n5928);
   U2760 : AOI222_X1 port map( A1 => n12, A2 => REGISTERS_82_8_port, B1 => n9, 
                           B2 => REGISTERS_84_8_port, C1 => n5, C2 => 
                           REGISTERS_83_8_port, ZN => n5937);
   U2761 : AOI222_X1 port map( A1 => n1143, A2 => REGISTERS_49_8_port, B1 => 
                           n1141, B2 => REGISTERS_51_8_port, C1 => n1138, C2 =>
                           REGISTERS_50_8_port, ZN => n4485);
   U2762 : AOI222_X1 port map( A1 => n725, A2 => REGISTERS_82_8_port, B1 => 
                           n723, B2 => REGISTERS_84_8_port, C1 => n720, C2 => 
                           REGISTERS_83_8_port, ZN => n4494);
   U2763 : AOI222_X1 port map( A1 => n79, A2 => REGISTERS_49_9_port, B1 => n77,
                           B2 => REGISTERS_51_9_port, C1 => n74, C2 => 
                           REGISTERS_50_9_port, ZN => n5887);
   U2764 : AOI222_X1 port map( A1 => n12, A2 => REGISTERS_82_9_port, B1 => n9, 
                           B2 => REGISTERS_84_9_port, C1 => n5, C2 => 
                           REGISTERS_83_9_port, ZN => n5896);
   U2765 : AOI222_X1 port map( A1 => n1143, A2 => REGISTERS_49_9_port, B1 => 
                           n1141, B2 => REGISTERS_51_9_port, C1 => n1138, C2 =>
                           REGISTERS_50_9_port, ZN => n4444);
   U2766 : AOI222_X1 port map( A1 => n725, A2 => REGISTERS_82_9_port, B1 => 
                           n723, B2 => REGISTERS_84_9_port, C1 => n720, C2 => 
                           REGISTERS_83_9_port, ZN => n4453);
   U2767 : AOI222_X1 port map( A1 => n79, A2 => REGISTERS_49_10_port, B1 => n77
                           , B2 => REGISTERS_51_10_port, C1 => n74, C2 => 
                           REGISTERS_50_10_port, ZN => n5846);
   U2768 : AOI222_X1 port map( A1 => n12, A2 => REGISTERS_82_10_port, B1 => n9,
                           B2 => REGISTERS_84_10_port, C1 => n5, C2 => 
                           REGISTERS_83_10_port, ZN => n5855);
   U2769 : AOI222_X1 port map( A1 => n1143, A2 => REGISTERS_49_10_port, B1 => 
                           n1141, B2 => REGISTERS_51_10_port, C1 => n1138, C2 
                           => REGISTERS_50_10_port, ZN => n4403);
   U2770 : AOI222_X1 port map( A1 => n725, A2 => REGISTERS_82_10_port, B1 => 
                           n723, B2 => REGISTERS_84_10_port, C1 => n720, C2 => 
                           REGISTERS_83_10_port, ZN => n4412);
   U2771 : AOI222_X1 port map( A1 => n79, A2 => REGISTERS_49_11_port, B1 => n77
                           , B2 => REGISTERS_51_11_port, C1 => n74, C2 => 
                           REGISTERS_50_11_port, ZN => n5805);
   U2772 : AOI222_X1 port map( A1 => n12, A2 => REGISTERS_82_11_port, B1 => n9,
                           B2 => REGISTERS_84_11_port, C1 => n5, C2 => 
                           REGISTERS_83_11_port, ZN => n5814);
   U2773 : AOI222_X1 port map( A1 => n1143, A2 => REGISTERS_49_11_port, B1 => 
                           n1141, B2 => REGISTERS_51_11_port, C1 => n1138, C2 
                           => REGISTERS_50_11_port, ZN => n4362);
   U2774 : AOI222_X1 port map( A1 => n725, A2 => REGISTERS_82_11_port, B1 => 
                           n723, B2 => REGISTERS_84_11_port, C1 => n720, C2 => 
                           REGISTERS_83_11_port, ZN => n4371);
   U2775 : AOI222_X1 port map( A1 => n432, A2 => REGISTERS_49_12_port, B1 => 
                           n77, B2 => REGISTERS_51_12_port, C1 => n74, C2 => 
                           REGISTERS_50_12_port, ZN => n5764);
   U2776 : AOI222_X1 port map( A1 => n13, A2 => REGISTERS_82_12_port, B1 => n9,
                           B2 => REGISTERS_84_12_port, C1 => n5, C2 => 
                           REGISTERS_83_12_port, ZN => n5773);
   U2777 : AOI222_X1 port map( A1 => n1144, A2 => REGISTERS_49_12_port, B1 => 
                           n1141, B2 => REGISTERS_51_12_port, C1 => n1138, C2 
                           => REGISTERS_50_12_port, ZN => n4321);
   U2778 : AOI222_X1 port map( A1 => n726, A2 => REGISTERS_82_12_port, B1 => 
                           n723, B2 => REGISTERS_84_12_port, C1 => n720, C2 => 
                           REGISTERS_83_12_port, ZN => n4330);
   U2779 : AOI222_X1 port map( A1 => n432, A2 => REGISTERS_49_13_port, B1 => 
                           n77, B2 => REGISTERS_51_13_port, C1 => n74, C2 => 
                           REGISTERS_50_13_port, ZN => n5723);
   U2780 : AOI222_X1 port map( A1 => n13, A2 => REGISTERS_82_13_port, B1 => n9,
                           B2 => REGISTERS_84_13_port, C1 => n5, C2 => 
                           REGISTERS_83_13_port, ZN => n5732);
   U2781 : AOI222_X1 port map( A1 => n1144, A2 => REGISTERS_49_13_port, B1 => 
                           n1141, B2 => REGISTERS_51_13_port, C1 => n1138, C2 
                           => REGISTERS_50_13_port, ZN => n4280);
   U2782 : AOI222_X1 port map( A1 => n726, A2 => REGISTERS_82_13_port, B1 => 
                           n723, B2 => REGISTERS_84_13_port, C1 => n720, C2 => 
                           REGISTERS_83_13_port, ZN => n4289);
   U2783 : AOI222_X1 port map( A1 => n432, A2 => REGISTERS_49_14_port, B1 => 
                           n77, B2 => REGISTERS_51_14_port, C1 => n74, C2 => 
                           REGISTERS_50_14_port, ZN => n5682);
   U2784 : AOI222_X1 port map( A1 => n13, A2 => REGISTERS_82_14_port, B1 => n9,
                           B2 => REGISTERS_84_14_port, C1 => n5, C2 => 
                           REGISTERS_83_14_port, ZN => n5691);
   U2785 : AOI222_X1 port map( A1 => n1144, A2 => REGISTERS_49_14_port, B1 => 
                           n1141, B2 => REGISTERS_51_14_port, C1 => n1138, C2 
                           => REGISTERS_50_14_port, ZN => n4239);
   U2786 : AOI222_X1 port map( A1 => n726, A2 => REGISTERS_82_14_port, B1 => 
                           n723, B2 => REGISTERS_84_14_port, C1 => n720, C2 => 
                           REGISTERS_83_14_port, ZN => n4248);
   U2787 : AOI222_X1 port map( A1 => n432, A2 => REGISTERS_49_15_port, B1 => 
                           n77, B2 => REGISTERS_51_15_port, C1 => n74, C2 => 
                           REGISTERS_50_15_port, ZN => n5641);
   U2788 : AOI222_X1 port map( A1 => n13, A2 => REGISTERS_82_15_port, B1 => n9,
                           B2 => REGISTERS_84_15_port, C1 => n5, C2 => 
                           REGISTERS_83_15_port, ZN => n5650);
   U2789 : AOI222_X1 port map( A1 => n1144, A2 => REGISTERS_49_15_port, B1 => 
                           n1141, B2 => REGISTERS_51_15_port, C1 => n1138, C2 
                           => REGISTERS_50_15_port, ZN => n4198);
   U2790 : AOI222_X1 port map( A1 => n726, A2 => REGISTERS_82_15_port, B1 => 
                           n723, B2 => REGISTERS_84_15_port, C1 => n720, C2 => 
                           REGISTERS_83_15_port, ZN => n4207);
   U2791 : AOI222_X1 port map( A1 => n432, A2 => REGISTERS_49_16_port, B1 => 
                           n77, B2 => REGISTERS_51_16_port, C1 => n74, C2 => 
                           REGISTERS_50_16_port, ZN => n5600);
   U2792 : AOI222_X1 port map( A1 => n13, A2 => REGISTERS_82_16_port, B1 => n9,
                           B2 => REGISTERS_84_16_port, C1 => n5, C2 => 
                           REGISTERS_83_16_port, ZN => n5609);
   U2793 : AOI222_X1 port map( A1 => n1144, A2 => REGISTERS_49_16_port, B1 => 
                           n1141, B2 => REGISTERS_51_16_port, C1 => n1138, C2 
                           => REGISTERS_50_16_port, ZN => n4157);
   U2794 : AOI222_X1 port map( A1 => n726, A2 => REGISTERS_82_16_port, B1 => 
                           n723, B2 => REGISTERS_84_16_port, C1 => n720, C2 => 
                           REGISTERS_83_16_port, ZN => n4166);
   U2795 : AOI222_X1 port map( A1 => n432, A2 => REGISTERS_49_17_port, B1 => 
                           n77, B2 => REGISTERS_51_17_port, C1 => n74, C2 => 
                           REGISTERS_50_17_port, ZN => n5559);
   U2796 : AOI222_X1 port map( A1 => n13, A2 => REGISTERS_82_17_port, B1 => n9,
                           B2 => REGISTERS_84_17_port, C1 => n5, C2 => 
                           REGISTERS_83_17_port, ZN => n5568);
   U2797 : AOI222_X1 port map( A1 => n1144, A2 => REGISTERS_49_17_port, B1 => 
                           n1141, B2 => REGISTERS_51_17_port, C1 => n1138, C2 
                           => REGISTERS_50_17_port, ZN => n4116);
   U2798 : AOI222_X1 port map( A1 => n726, A2 => REGISTERS_82_17_port, B1 => 
                           n723, B2 => REGISTERS_84_17_port, C1 => n720, C2 => 
                           REGISTERS_83_17_port, ZN => n4125);
   U2799 : AOI222_X1 port map( A1 => n432, A2 => REGISTERS_49_18_port, B1 => 
                           n77, B2 => REGISTERS_51_18_port, C1 => n74, C2 => 
                           REGISTERS_50_18_port, ZN => n5518);
   U2800 : AOI222_X1 port map( A1 => n13, A2 => REGISTERS_82_18_port, B1 => n9,
                           B2 => REGISTERS_84_18_port, C1 => n5, C2 => 
                           REGISTERS_83_18_port, ZN => n5527);
   U2801 : AOI222_X1 port map( A1 => n1144, A2 => REGISTERS_49_18_port, B1 => 
                           n1141, B2 => REGISTERS_51_18_port, C1 => n1138, C2 
                           => REGISTERS_50_18_port, ZN => n4075);
   U2802 : AOI222_X1 port map( A1 => n726, A2 => REGISTERS_82_18_port, B1 => 
                           n723, B2 => REGISTERS_84_18_port, C1 => n720, C2 => 
                           REGISTERS_83_18_port, ZN => n4084);
   U2803 : AOI222_X1 port map( A1 => n432, A2 => REGISTERS_49_19_port, B1 => 
                           n77, B2 => REGISTERS_51_19_port, C1 => n74, C2 => 
                           REGISTERS_50_19_port, ZN => n5477);
   U2804 : AOI222_X1 port map( A1 => n13, A2 => REGISTERS_82_19_port, B1 => n9,
                           B2 => REGISTERS_84_19_port, C1 => n5, C2 => 
                           REGISTERS_83_19_port, ZN => n5486);
   U2805 : AOI222_X1 port map( A1 => n1144, A2 => REGISTERS_49_19_port, B1 => 
                           n1141, B2 => REGISTERS_51_19_port, C1 => n1138, C2 
                           => REGISTERS_50_19_port, ZN => n4034);
   U2806 : AOI222_X1 port map( A1 => n726, A2 => REGISTERS_82_19_port, B1 => 
                           n723, B2 => REGISTERS_84_19_port, C1 => n720, C2 => 
                           REGISTERS_83_19_port, ZN => n4043);
   U2807 : AOI222_X1 port map( A1 => n432, A2 => REGISTERS_49_20_port, B1 => 
                           n76, B2 => REGISTERS_51_20_port, C1 => n73, C2 => 
                           REGISTERS_50_20_port, ZN => n5436);
   U2808 : AOI222_X1 port map( A1 => n13, A2 => REGISTERS_82_20_port, B1 => n8,
                           B2 => REGISTERS_84_20_port, C1 => n4, C2 => 
                           REGISTERS_83_20_port, ZN => n5445);
   U2809 : AOI222_X1 port map( A1 => n1144, A2 => REGISTERS_49_20_port, B1 => 
                           n1140, B2 => REGISTERS_51_20_port, C1 => n1137, C2 
                           => REGISTERS_50_20_port, ZN => n3993);
   U2810 : AOI222_X1 port map( A1 => n726, A2 => REGISTERS_82_20_port, B1 => 
                           n722, B2 => REGISTERS_84_20_port, C1 => n719, C2 => 
                           REGISTERS_83_20_port, ZN => n4002);
   U2811 : AOI222_X1 port map( A1 => n432, A2 => REGISTERS_49_21_port, B1 => 
                           n76, B2 => REGISTERS_51_21_port, C1 => n73, C2 => 
                           REGISTERS_50_21_port, ZN => n5395);
   U2812 : AOI222_X1 port map( A1 => n13, A2 => REGISTERS_82_21_port, B1 => n8,
                           B2 => REGISTERS_84_21_port, C1 => n4, C2 => 
                           REGISTERS_83_21_port, ZN => n5404);
   U2813 : AOI222_X1 port map( A1 => n1144, A2 => REGISTERS_49_21_port, B1 => 
                           n1140, B2 => REGISTERS_51_21_port, C1 => n1137, C2 
                           => REGISTERS_50_21_port, ZN => n3952);
   U2814 : AOI222_X1 port map( A1 => n726, A2 => REGISTERS_82_21_port, B1 => 
                           n722, B2 => REGISTERS_84_21_port, C1 => n719, C2 => 
                           REGISTERS_83_21_port, ZN => n3961);
   U2815 : AOI222_X1 port map( A1 => n432, A2 => REGISTERS_49_22_port, B1 => 
                           n76, B2 => REGISTERS_51_22_port, C1 => n73, C2 => 
                           REGISTERS_50_22_port, ZN => n5354);
   U2816 : AOI222_X1 port map( A1 => n13, A2 => REGISTERS_82_22_port, B1 => n8,
                           B2 => REGISTERS_84_22_port, C1 => n4, C2 => 
                           REGISTERS_83_22_port, ZN => n5363);
   U2817 : AOI222_X1 port map( A1 => n1144, A2 => REGISTERS_49_22_port, B1 => 
                           n1140, B2 => REGISTERS_51_22_port, C1 => n1137, C2 
                           => REGISTERS_50_22_port, ZN => n3911);
   U2818 : AOI222_X1 port map( A1 => n726, A2 => REGISTERS_82_22_port, B1 => 
                           n722, B2 => REGISTERS_84_22_port, C1 => n719, C2 => 
                           REGISTERS_83_22_port, ZN => n3920);
   U2819 : AOI222_X1 port map( A1 => n432, A2 => REGISTERS_49_23_port, B1 => 
                           n76, B2 => REGISTERS_51_23_port, C1 => n73, C2 => 
                           REGISTERS_50_23_port, ZN => n5313);
   U2820 : AOI222_X1 port map( A1 => n13, A2 => REGISTERS_82_23_port, B1 => n8,
                           B2 => REGISTERS_84_23_port, C1 => n4, C2 => 
                           REGISTERS_83_23_port, ZN => n5322);
   U2821 : AOI222_X1 port map( A1 => n1144, A2 => REGISTERS_49_23_port, B1 => 
                           n1140, B2 => REGISTERS_51_23_port, C1 => n1137, C2 
                           => REGISTERS_50_23_port, ZN => n3870);
   U2822 : AOI222_X1 port map( A1 => n726, A2 => REGISTERS_82_23_port, B1 => 
                           n722, B2 => REGISTERS_84_23_port, C1 => n719, C2 => 
                           REGISTERS_83_23_port, ZN => n3879);
   U2823 : AOI222_X1 port map( A1 => n433, A2 => REGISTERS_49_24_port, B1 => 
                           n76, B2 => REGISTERS_51_24_port, C1 => n73, C2 => 
                           REGISTERS_50_24_port, ZN => n5272);
   U2824 : AOI222_X1 port map( A1 => n14, A2 => REGISTERS_82_24_port, B1 => n8,
                           B2 => REGISTERS_84_24_port, C1 => n4, C2 => 
                           REGISTERS_83_24_port, ZN => n5281);
   U2825 : AOI222_X1 port map( A1 => n1145, A2 => REGISTERS_49_24_port, B1 => 
                           n1140, B2 => REGISTERS_51_24_port, C1 => n1137, C2 
                           => REGISTERS_50_24_port, ZN => n3829);
   U2826 : AOI222_X1 port map( A1 => n727, A2 => REGISTERS_82_24_port, B1 => 
                           n722, B2 => REGISTERS_84_24_port, C1 => n719, C2 => 
                           REGISTERS_83_24_port, ZN => n3838);
   U2827 : AOI222_X1 port map( A1 => n433, A2 => REGISTERS_49_25_port, B1 => 
                           n76, B2 => REGISTERS_51_25_port, C1 => n73, C2 => 
                           REGISTERS_50_25_port, ZN => n5231);
   U2828 : AOI222_X1 port map( A1 => n14, A2 => REGISTERS_82_25_port, B1 => n8,
                           B2 => REGISTERS_84_25_port, C1 => n4, C2 => 
                           REGISTERS_83_25_port, ZN => n5240);
   U2829 : AOI222_X1 port map( A1 => n1145, A2 => REGISTERS_49_25_port, B1 => 
                           n1140, B2 => REGISTERS_51_25_port, C1 => n1137, C2 
                           => REGISTERS_50_25_port, ZN => n3788);
   U2830 : AOI222_X1 port map( A1 => n727, A2 => REGISTERS_82_25_port, B1 => 
                           n722, B2 => REGISTERS_84_25_port, C1 => n719, C2 => 
                           REGISTERS_83_25_port, ZN => n3797);
   U2831 : AOI222_X1 port map( A1 => n433, A2 => REGISTERS_49_26_port, B1 => 
                           n76, B2 => REGISTERS_51_26_port, C1 => n73, C2 => 
                           REGISTERS_50_26_port, ZN => n5190);
   U2832 : AOI222_X1 port map( A1 => n14, A2 => REGISTERS_82_26_port, B1 => n8,
                           B2 => REGISTERS_84_26_port, C1 => n4, C2 => 
                           REGISTERS_83_26_port, ZN => n5199);
   U2833 : AOI222_X1 port map( A1 => n1145, A2 => REGISTERS_49_26_port, B1 => 
                           n1140, B2 => REGISTERS_51_26_port, C1 => n1137, C2 
                           => REGISTERS_50_26_port, ZN => n3747);
   U2834 : AOI222_X1 port map( A1 => n727, A2 => REGISTERS_82_26_port, B1 => 
                           n722, B2 => REGISTERS_84_26_port, C1 => n719, C2 => 
                           REGISTERS_83_26_port, ZN => n3756);
   U2835 : AOI222_X1 port map( A1 => n433, A2 => REGISTERS_49_27_port, B1 => 
                           n76, B2 => REGISTERS_51_27_port, C1 => n73, C2 => 
                           REGISTERS_50_27_port, ZN => n5149);
   U2836 : AOI222_X1 port map( A1 => n14, A2 => REGISTERS_82_27_port, B1 => n8,
                           B2 => REGISTERS_84_27_port, C1 => n4, C2 => 
                           REGISTERS_83_27_port, ZN => n5158);
   U2837 : AOI222_X1 port map( A1 => n1145, A2 => REGISTERS_49_27_port, B1 => 
                           n1140, B2 => REGISTERS_51_27_port, C1 => n1137, C2 
                           => REGISTERS_50_27_port, ZN => n3706);
   U2838 : AOI222_X1 port map( A1 => n727, A2 => REGISTERS_82_27_port, B1 => 
                           n722, B2 => REGISTERS_84_27_port, C1 => n719, C2 => 
                           REGISTERS_83_27_port, ZN => n3715);
   U2839 : AOI222_X1 port map( A1 => n433, A2 => REGISTERS_49_28_port, B1 => 
                           n76, B2 => REGISTERS_51_28_port, C1 => n73, C2 => 
                           REGISTERS_50_28_port, ZN => n5108);
   U2840 : AOI222_X1 port map( A1 => n14, A2 => REGISTERS_82_28_port, B1 => n8,
                           B2 => REGISTERS_84_28_port, C1 => n4, C2 => 
                           REGISTERS_83_28_port, ZN => n5117);
   U2841 : AOI222_X1 port map( A1 => n1145, A2 => REGISTERS_49_28_port, B1 => 
                           n1140, B2 => REGISTERS_51_28_port, C1 => n1137, C2 
                           => REGISTERS_50_28_port, ZN => n3665);
   U2842 : AOI222_X1 port map( A1 => n727, A2 => REGISTERS_82_28_port, B1 => 
                           n722, B2 => REGISTERS_84_28_port, C1 => n719, C2 => 
                           REGISTERS_83_28_port, ZN => n3674);
   U2843 : AOI222_X1 port map( A1 => n433, A2 => REGISTERS_49_29_port, B1 => 
                           n76, B2 => REGISTERS_51_29_port, C1 => n73, C2 => 
                           REGISTERS_50_29_port, ZN => n5067);
   U2844 : AOI222_X1 port map( A1 => n14, A2 => REGISTERS_82_29_port, B1 => n8,
                           B2 => REGISTERS_84_29_port, C1 => n4, C2 => 
                           REGISTERS_83_29_port, ZN => n5076);
   U2845 : AOI222_X1 port map( A1 => n1145, A2 => REGISTERS_49_29_port, B1 => 
                           n1140, B2 => REGISTERS_51_29_port, C1 => n1137, C2 
                           => REGISTERS_50_29_port, ZN => n3624);
   U2846 : AOI222_X1 port map( A1 => n727, A2 => REGISTERS_82_29_port, B1 => 
                           n722, B2 => REGISTERS_84_29_port, C1 => n719, C2 => 
                           REGISTERS_83_29_port, ZN => n3633);
   U2847 : AOI222_X1 port map( A1 => n433, A2 => REGISTERS_49_30_port, B1 => 
                           n76, B2 => REGISTERS_51_30_port, C1 => n73, C2 => 
                           REGISTERS_50_30_port, ZN => n5026);
   U2848 : AOI222_X1 port map( A1 => n14, A2 => REGISTERS_82_30_port, B1 => n8,
                           B2 => REGISTERS_84_30_port, C1 => n4, C2 => 
                           REGISTERS_83_30_port, ZN => n5035);
   U2849 : AOI222_X1 port map( A1 => n1145, A2 => REGISTERS_49_30_port, B1 => 
                           n1140, B2 => REGISTERS_51_30_port, C1 => n1137, C2 
                           => REGISTERS_50_30_port, ZN => n3583);
   U2850 : AOI222_X1 port map( A1 => n727, A2 => REGISTERS_82_30_port, B1 => 
                           n722, B2 => REGISTERS_84_30_port, C1 => n719, C2 => 
                           REGISTERS_83_30_port, ZN => n3592);
   U2851 : AOI222_X1 port map( A1 => n433, A2 => REGISTERS_49_31_port, B1 => 
                           n76, B2 => REGISTERS_51_31_port, C1 => n73, C2 => 
                           REGISTERS_50_31_port, ZN => n4941);
   U2852 : AOI222_X1 port map( A1 => n14, A2 => REGISTERS_82_31_port, B1 => n8,
                           B2 => REGISTERS_84_31_port, C1 => n4, C2 => 
                           REGISTERS_83_31_port, ZN => n4972);
   U2853 : AOI222_X1 port map( A1 => n1145, A2 => REGISTERS_49_31_port, B1 => 
                           n1140, B2 => REGISTERS_51_31_port, C1 => n1137, C2 
                           => REGISTERS_50_31_port, ZN => n3498);
   U2854 : AOI222_X1 port map( A1 => n727, A2 => REGISTERS_82_31_port, B1 => 
                           n722, B2 => REGISTERS_84_31_port, C1 => n719, C2 => 
                           REGISTERS_83_31_port, ZN => n3529);
   U2855 : NOR4_X1 port map( A1 => n6292, A2 => n6293, A3 => n6294, A4 => n6295
                           , ZN => n6291);
   U2856 : OAI22_X1 port map( A1 => n1871, A2 => n488, B1 => n1903, B2 => n485,
                           ZN => n6295);
   U2857 : OAI222_X1 port map( A1 => n2159_port, A2 => n464, B1 => n2191, B2 =>
                           n461, C1 => n2127, C2 => n458, ZN => n6292);
   U2858 : OAI222_X1 port map( A1 => n2063, A2 => n473, B1 => n2095, B2 => n470
                           , C1 => n2031, C2 => n467, ZN => n6293);
   U2859 : NOR4_X1 port map( A1 => n6305, A2 => n6306, A3 => n6307, A4 => n6308
                           , ZN => n6304);
   U2860 : OAI22_X1 port map( A1 => n2223, A2 => n70, B1 => n2255, B2 => n67, 
                           ZN => n6308);
   U2861 : OAI222_X1 port map( A1 => n2511, A2 => n46, B1 => n2543, B2 => n43, 
                           C1 => n2479, C2 => n40, ZN => n6305);
   U2862 : OAI222_X1 port map( A1 => n2415, A2 => n55, B1 => n2447, B2 => n52, 
                           C1 => n2383, C2 => n49, ZN => n6306);
   U2863 : NOR4_X1 port map( A1 => n4849, A2 => n4850, A3 => n4851, A4 => n4852
                           , ZN => n4848);
   U2864 : OAI22_X1 port map( A1 => n1871, A2 => n1296, B1 => n1903, B2 => 
                           n1197, ZN => n4852);
   U2865 : OAI222_X1 port map( A1 => n2159_port, A2 => n1176, B1 => n2191, B2 
                           => n1173, C1 => n2127, C2 => n1170, ZN => n4849);
   U2866 : OAI222_X1 port map( A1 => n2063, A2 => n1185, B1 => n2095, B2 => 
                           n1182, C1 => n2031, C2 => n1179, ZN => n4850);
   U2867 : NOR4_X1 port map( A1 => n4862, A2 => n4863, A3 => n4864, A4 => n4865
                           , ZN => n4861);
   U2868 : OAI22_X1 port map( A1 => n2223, A2 => n782, B1 => n2255, B2 => n779,
                           ZN => n4865);
   U2869 : OAI222_X1 port map( A1 => n2511, A2 => n758, B1 => n2543, B2 => n755
                           , C1 => n2479, C2 => n752, ZN => n4862);
   U2870 : OAI222_X1 port map( A1 => n2415, A2 => n767, B1 => n2447, B2 => n764
                           , C1 => n2383, C2 => n761, ZN => n4863);
   U2871 : NOR4_X1 port map( A1 => n6219, A2 => n6220, A3 => n6221, A4 => n6222
                           , ZN => n6218);
   U2872 : OAI22_X1 port map( A1 => n1870, A2 => n488, B1 => n1902, B2 => n485,
                           ZN => n6222);
   U2873 : OAI222_X1 port map( A1 => n2158_port, A2 => n464, B1 => n2190, B2 =>
                           n461, C1 => n2126, C2 => n458, ZN => n6219);
   U2874 : OAI222_X1 port map( A1 => n2062, A2 => n473, B1 => n2094, B2 => n470
                           , C1 => n2030, C2 => n467, ZN => n6220);
   U2875 : NOR4_X1 port map( A1 => n6228, A2 => n6229, A3 => n6230, A4 => n6231
                           , ZN => n6227);
   U2876 : OAI22_X1 port map( A1 => n2222, A2 => n70, B1 => n2254, B2 => n67, 
                           ZN => n6231);
   U2877 : OAI222_X1 port map( A1 => n2510, A2 => n46, B1 => n2542, B2 => n43, 
                           C1 => n2478, C2 => n40, ZN => n6228);
   U2878 : OAI222_X1 port map( A1 => n2414, A2 => n55, B1 => n2446, B2 => n52, 
                           C1 => n2382, C2 => n49, ZN => n6229);
   U2879 : NOR4_X1 port map( A1 => n4776, A2 => n4777, A3 => n4778, A4 => n4779
                           , ZN => n4775);
   U2880 : OAI22_X1 port map( A1 => n1870, A2 => n1296, B1 => n1902, B2 => 
                           n1197, ZN => n4779);
   U2881 : OAI222_X1 port map( A1 => n2158_port, A2 => n1176, B1 => n2190, B2 
                           => n1173, C1 => n2126, C2 => n1170, ZN => n4776);
   U2882 : OAI222_X1 port map( A1 => n2062, A2 => n1185, B1 => n2094, B2 => 
                           n1182, C1 => n2030, C2 => n1179, ZN => n4777);
   U2883 : NOR4_X1 port map( A1 => n4785, A2 => n4786, A3 => n4787, A4 => n4788
                           , ZN => n4784);
   U2884 : OAI22_X1 port map( A1 => n2222, A2 => n782, B1 => n2254, B2 => n779,
                           ZN => n4788);
   U2885 : OAI222_X1 port map( A1 => n2510, A2 => n758, B1 => n2542, B2 => n755
                           , C1 => n2478, C2 => n752, ZN => n4785);
   U2886 : OAI222_X1 port map( A1 => n2414, A2 => n767, B1 => n2446, B2 => n764
                           , C1 => n2382, C2 => n761, ZN => n4786);
   U2887 : NOR4_X1 port map( A1 => n6178, A2 => n6179, A3 => n6180, A4 => n6181
                           , ZN => n6177);
   U2888 : OAI22_X1 port map( A1 => n1869, A2 => n488, B1 => n1901, B2 => n485,
                           ZN => n6181);
   U2889 : OAI222_X1 port map( A1 => n2157_port, A2 => n464, B1 => n2189, B2 =>
                           n461, C1 => n2125, C2 => n458, ZN => n6178);
   U2890 : OAI222_X1 port map( A1 => n2061, A2 => n473, B1 => n2093, B2 => n470
                           , C1 => n2029, C2 => n467, ZN => n6179);
   U2891 : NOR4_X1 port map( A1 => n6187, A2 => n6188, A3 => n6189, A4 => n6190
                           , ZN => n6186);
   U2892 : OAI22_X1 port map( A1 => n2221, A2 => n70, B1 => n2253, B2 => n67, 
                           ZN => n6190);
   U2893 : OAI222_X1 port map( A1 => n2509, A2 => n46, B1 => n2541, B2 => n43, 
                           C1 => n2477, C2 => n40, ZN => n6187);
   U2894 : OAI222_X1 port map( A1 => n2413, A2 => n55, B1 => n2445, B2 => n52, 
                           C1 => n2381, C2 => n49, ZN => n6188);
   U2895 : NOR4_X1 port map( A1 => n4735, A2 => n4736, A3 => n4737, A4 => n4738
                           , ZN => n4734);
   U2896 : OAI22_X1 port map( A1 => n1869, A2 => n1296, B1 => n1901, B2 => 
                           n1197, ZN => n4738);
   U2897 : OAI222_X1 port map( A1 => n2157_port, A2 => n1176, B1 => n2189, B2 
                           => n1173, C1 => n2125, C2 => n1170, ZN => n4735);
   U2898 : OAI222_X1 port map( A1 => n2061, A2 => n1185, B1 => n2093, B2 => 
                           n1182, C1 => n2029, C2 => n1179, ZN => n4736);
   U2899 : NOR4_X1 port map( A1 => n4744, A2 => n4745, A3 => n4746, A4 => n4747
                           , ZN => n4743);
   U2900 : OAI22_X1 port map( A1 => n2221, A2 => n782, B1 => n2253, B2 => n779,
                           ZN => n4747);
   U2901 : OAI222_X1 port map( A1 => n2509, A2 => n758, B1 => n2541, B2 => n755
                           , C1 => n2477, C2 => n752, ZN => n4744);
   U2902 : OAI222_X1 port map( A1 => n2413, A2 => n767, B1 => n2445, B2 => n764
                           , C1 => n2381, C2 => n761, ZN => n4745);
   U2903 : NOR4_X1 port map( A1 => n6137, A2 => n6138, A3 => n6139, A4 => n6140
                           , ZN => n6136);
   U2904 : OAI22_X1 port map( A1 => n1868, A2 => n488, B1 => n1900, B2 => n485,
                           ZN => n6140);
   U2905 : OAI222_X1 port map( A1 => n2156_port, A2 => n464, B1 => n2188, B2 =>
                           n461, C1 => n2124, C2 => n458, ZN => n6137);
   U2906 : OAI222_X1 port map( A1 => n2060, A2 => n473, B1 => n2092, B2 => n470
                           , C1 => n2028, C2 => n467, ZN => n6138);
   U2907 : NOR4_X1 port map( A1 => n6146, A2 => n6147, A3 => n6148, A4 => n6149
                           , ZN => n6145);
   U2908 : OAI22_X1 port map( A1 => n2220, A2 => n70, B1 => n2252, B2 => n67, 
                           ZN => n6149);
   U2909 : OAI222_X1 port map( A1 => n2508, A2 => n46, B1 => n2540, B2 => n43, 
                           C1 => n2476, C2 => n40, ZN => n6146);
   U2910 : OAI222_X1 port map( A1 => n2412, A2 => n55, B1 => n2444, B2 => n52, 
                           C1 => n2380, C2 => n49, ZN => n6147);
   U2911 : NOR4_X1 port map( A1 => n4694, A2 => n4695, A3 => n4696, A4 => n4697
                           , ZN => n4693);
   U2912 : OAI22_X1 port map( A1 => n1868, A2 => n1296, B1 => n1900, B2 => 
                           n1197, ZN => n4697);
   U2913 : OAI222_X1 port map( A1 => n2156_port, A2 => n1176, B1 => n2188, B2 
                           => n1173, C1 => n2124, C2 => n1170, ZN => n4694);
   U2914 : OAI222_X1 port map( A1 => n2060, A2 => n1185, B1 => n2092, B2 => 
                           n1182, C1 => n2028, C2 => n1179, ZN => n4695);
   U2915 : NOR4_X1 port map( A1 => n4703, A2 => n4704, A3 => n4705, A4 => n4706
                           , ZN => n4702);
   U2916 : OAI22_X1 port map( A1 => n2220, A2 => n782, B1 => n2252, B2 => n779,
                           ZN => n4706);
   U2917 : OAI222_X1 port map( A1 => n2508, A2 => n758, B1 => n2540, B2 => n755
                           , C1 => n2476, C2 => n752, ZN => n4703);
   U2918 : OAI222_X1 port map( A1 => n2412, A2 => n767, B1 => n2444, B2 => n764
                           , C1 => n2380, C2 => n761, ZN => n4704);
   U2919 : NOR4_X1 port map( A1 => n6096, A2 => n6097, A3 => n6098, A4 => n6099
                           , ZN => n6095);
   U2920 : OAI22_X1 port map( A1 => n1867, A2 => n488, B1 => n1899, B2 => n485,
                           ZN => n6099);
   U2921 : OAI222_X1 port map( A1 => n2155_port, A2 => n464, B1 => n2187, B2 =>
                           n461, C1 => n2123, C2 => n458, ZN => n6096);
   U2922 : OAI222_X1 port map( A1 => n2059, A2 => n473, B1 => n2091, B2 => n470
                           , C1 => n2027, C2 => n467, ZN => n6097);
   U2923 : NOR4_X1 port map( A1 => n6105, A2 => n6106, A3 => n6107, A4 => n6108
                           , ZN => n6104);
   U2924 : OAI22_X1 port map( A1 => n2219, A2 => n70, B1 => n2251, B2 => n67, 
                           ZN => n6108);
   U2925 : OAI222_X1 port map( A1 => n2507, A2 => n46, B1 => n2539, B2 => n43, 
                           C1 => n2475, C2 => n40, ZN => n6105);
   U2926 : OAI222_X1 port map( A1 => n2411, A2 => n55, B1 => n2443, B2 => n52, 
                           C1 => n2379, C2 => n49, ZN => n6106);
   U2927 : NOR4_X1 port map( A1 => n4653, A2 => n4654, A3 => n4655, A4 => n4656
                           , ZN => n4652);
   U2928 : OAI22_X1 port map( A1 => n1867, A2 => n1296, B1 => n1899, B2 => 
                           n1197, ZN => n4656);
   U2929 : OAI222_X1 port map( A1 => n2155_port, A2 => n1176, B1 => n2187, B2 
                           => n1173, C1 => n2123, C2 => n1170, ZN => n4653);
   U2930 : OAI222_X1 port map( A1 => n2059, A2 => n1185, B1 => n2091, B2 => 
                           n1182, C1 => n2027, C2 => n1179, ZN => n4654);
   U2931 : NOR4_X1 port map( A1 => n4662, A2 => n4663, A3 => n4664, A4 => n4665
                           , ZN => n4661);
   U2932 : OAI22_X1 port map( A1 => n2219, A2 => n782, B1 => n2251, B2 => n779,
                           ZN => n4665);
   U2933 : OAI222_X1 port map( A1 => n2507, A2 => n758, B1 => n2539, B2 => n755
                           , C1 => n2475, C2 => n752, ZN => n4662);
   U2934 : OAI222_X1 port map( A1 => n2411, A2 => n767, B1 => n2443, B2 => n764
                           , C1 => n2379, C2 => n761, ZN => n4663);
   U2935 : NOR4_X1 port map( A1 => n6055, A2 => n6056, A3 => n6057, A4 => n6058
                           , ZN => n6054);
   U2936 : OAI22_X1 port map( A1 => n1866, A2 => n488, B1 => n1898, B2 => n485,
                           ZN => n6058);
   U2937 : OAI222_X1 port map( A1 => n2154_port, A2 => n464, B1 => n2186, B2 =>
                           n461, C1 => n2122, C2 => n458, ZN => n6055);
   U2938 : OAI222_X1 port map( A1 => n2058, A2 => n473, B1 => n2090, B2 => n470
                           , C1 => n2026, C2 => n467, ZN => n6056);
   U2939 : NOR4_X1 port map( A1 => n6064, A2 => n6065, A3 => n6066, A4 => n6067
                           , ZN => n6063);
   U2940 : OAI22_X1 port map( A1 => n2218, A2 => n70, B1 => n2250, B2 => n67, 
                           ZN => n6067);
   U2941 : OAI222_X1 port map( A1 => n2506, A2 => n46, B1 => n2538, B2 => n43, 
                           C1 => n2474, C2 => n40, ZN => n6064);
   U2942 : OAI222_X1 port map( A1 => n2410, A2 => n55, B1 => n2442, B2 => n52, 
                           C1 => n2378, C2 => n49, ZN => n6065);
   U2943 : NOR4_X1 port map( A1 => n4612, A2 => n4613, A3 => n4614, A4 => n4615
                           , ZN => n4611);
   U2944 : OAI22_X1 port map( A1 => n1866, A2 => n1296, B1 => n1898, B2 => 
                           n1197, ZN => n4615);
   U2945 : OAI222_X1 port map( A1 => n2154_port, A2 => n1176, B1 => n2186, B2 
                           => n1173, C1 => n2122, C2 => n1170, ZN => n4612);
   U2946 : OAI222_X1 port map( A1 => n2058, A2 => n1185, B1 => n2090, B2 => 
                           n1182, C1 => n2026, C2 => n1179, ZN => n4613);
   U2947 : NOR4_X1 port map( A1 => n4621, A2 => n4622, A3 => n4623, A4 => n4624
                           , ZN => n4620);
   U2948 : OAI22_X1 port map( A1 => n2218, A2 => n782, B1 => n2250, B2 => n779,
                           ZN => n4624);
   U2949 : OAI222_X1 port map( A1 => n2506, A2 => n758, B1 => n2538, B2 => n755
                           , C1 => n2474, C2 => n752, ZN => n4621);
   U2950 : OAI222_X1 port map( A1 => n2410, A2 => n767, B1 => n2442, B2 => n764
                           , C1 => n2378, C2 => n761, ZN => n4622);
   U2951 : NOR4_X1 port map( A1 => n6014, A2 => n6015, A3 => n6016, A4 => n6017
                           , ZN => n6013);
   U2952 : OAI22_X1 port map( A1 => n1865, A2 => n488, B1 => n1897, B2 => n485,
                           ZN => n6017);
   U2953 : OAI222_X1 port map( A1 => n2153_port, A2 => n464, B1 => n2185, B2 =>
                           n461, C1 => n2121, C2 => n458, ZN => n6014);
   U2954 : OAI222_X1 port map( A1 => n2057, A2 => n473, B1 => n2089, B2 => n470
                           , C1 => n2025, C2 => n467, ZN => n6015);
   U2955 : NOR4_X1 port map( A1 => n6023, A2 => n6024, A3 => n6025, A4 => n6026
                           , ZN => n6022);
   U2956 : OAI22_X1 port map( A1 => n2217, A2 => n70, B1 => n2249, B2 => n67, 
                           ZN => n6026);
   U2957 : OAI222_X1 port map( A1 => n2505, A2 => n46, B1 => n2537, B2 => n43, 
                           C1 => n2473, C2 => n40, ZN => n6023);
   U2958 : OAI222_X1 port map( A1 => n2409, A2 => n55, B1 => n2441, B2 => n52, 
                           C1 => n2377, C2 => n49, ZN => n6024);
   U2959 : NOR4_X1 port map( A1 => n4571, A2 => n4572, A3 => n4573, A4 => n4574
                           , ZN => n4570);
   U2960 : OAI22_X1 port map( A1 => n1865, A2 => n1296, B1 => n1897, B2 => 
                           n1197, ZN => n4574);
   U2961 : OAI222_X1 port map( A1 => n2153_port, A2 => n1176, B1 => n2185, B2 
                           => n1173, C1 => n2121, C2 => n1170, ZN => n4571);
   U2962 : OAI222_X1 port map( A1 => n2057, A2 => n1185, B1 => n2089, B2 => 
                           n1182, C1 => n2025, C2 => n1179, ZN => n4572);
   U2963 : NOR4_X1 port map( A1 => n4580, A2 => n4581, A3 => n4582, A4 => n4583
                           , ZN => n4579);
   U2964 : OAI22_X1 port map( A1 => n2217, A2 => n782, B1 => n2249, B2 => n779,
                           ZN => n4583);
   U2965 : OAI222_X1 port map( A1 => n2505, A2 => n758, B1 => n2537, B2 => n755
                           , C1 => n2473, C2 => n752, ZN => n4580);
   U2966 : OAI222_X1 port map( A1 => n2409, A2 => n767, B1 => n2441, B2 => n764
                           , C1 => n2377, C2 => n761, ZN => n4581);
   U2967 : NOR4_X1 port map( A1 => n5973, A2 => n5974, A3 => n5975, A4 => n5976
                           , ZN => n5972);
   U2968 : OAI22_X1 port map( A1 => n1864, A2 => n488, B1 => n1896, B2 => n485,
                           ZN => n5976);
   U2969 : OAI222_X1 port map( A1 => n2152, A2 => n464, B1 => n2184, B2 => n461
                           , C1 => n2120, C2 => n458, ZN => n5973);
   U2970 : OAI222_X1 port map( A1 => n2056, A2 => n473, B1 => n2088, B2 => n470
                           , C1 => n2024, C2 => n467, ZN => n5974);
   U2971 : NOR4_X1 port map( A1 => n5982, A2 => n5983, A3 => n5984, A4 => n5985
                           , ZN => n5981);
   U2972 : OAI22_X1 port map( A1 => n2216, A2 => n70, B1 => n2248, B2 => n67, 
                           ZN => n5985);
   U2973 : OAI222_X1 port map( A1 => n2504, A2 => n46, B1 => n2536, B2 => n43, 
                           C1 => n2472, C2 => n40, ZN => n5982);
   U2974 : OAI222_X1 port map( A1 => n2408, A2 => n55, B1 => n2440, B2 => n52, 
                           C1 => n2376, C2 => n49, ZN => n5983);
   U2975 : NOR4_X1 port map( A1 => n4530, A2 => n4531, A3 => n4532, A4 => n4533
                           , ZN => n4529);
   U2976 : OAI22_X1 port map( A1 => n1864, A2 => n1296, B1 => n1896, B2 => 
                           n1197, ZN => n4533);
   U2977 : OAI222_X1 port map( A1 => n2152, A2 => n1176, B1 => n2184, B2 => 
                           n1173, C1 => n2120, C2 => n1170, ZN => n4530);
   U2978 : OAI222_X1 port map( A1 => n2056, A2 => n1185, B1 => n2088, B2 => 
                           n1182, C1 => n2024, C2 => n1179, ZN => n4531);
   U2979 : NOR4_X1 port map( A1 => n4539, A2 => n4540, A3 => n4541, A4 => n4542
                           , ZN => n4538);
   U2980 : OAI22_X1 port map( A1 => n2216, A2 => n782, B1 => n2248, B2 => n779,
                           ZN => n4542);
   U2981 : OAI222_X1 port map( A1 => n2504, A2 => n758, B1 => n2536, B2 => n755
                           , C1 => n2472, C2 => n752, ZN => n4539);
   U2982 : OAI222_X1 port map( A1 => n2408, A2 => n767, B1 => n2440, B2 => n764
                           , C1 => n2376, C2 => n761, ZN => n4540);
   U2983 : NOR4_X1 port map( A1 => n5932, A2 => n5933, A3 => n5934, A4 => n5935
                           , ZN => n5931);
   U2984 : OAI22_X1 port map( A1 => n1863, A2 => n488, B1 => n1895, B2 => n485,
                           ZN => n5935);
   U2985 : OAI222_X1 port map( A1 => n2151_port, A2 => n464, B1 => n2183, B2 =>
                           n461, C1 => n2119, C2 => n458, ZN => n5932);
   U2986 : OAI222_X1 port map( A1 => n2055, A2 => n473, B1 => n2087, B2 => n470
                           , C1 => n2023, C2 => n467, ZN => n5933);
   U2987 : NOR4_X1 port map( A1 => n5941, A2 => n5942, A3 => n5943, A4 => n5944
                           , ZN => n5940);
   U2988 : OAI22_X1 port map( A1 => n2215, A2 => n70, B1 => n2247, B2 => n67, 
                           ZN => n5944);
   U2989 : OAI222_X1 port map( A1 => n2503, A2 => n46, B1 => n2535, B2 => n43, 
                           C1 => n2471, C2 => n40, ZN => n5941);
   U2990 : OAI222_X1 port map( A1 => n2407, A2 => n55, B1 => n2439, B2 => n52, 
                           C1 => n2375, C2 => n49, ZN => n5942);
   U2991 : NOR4_X1 port map( A1 => n4489, A2 => n4490, A3 => n4491, A4 => n4492
                           , ZN => n4488);
   U2992 : OAI22_X1 port map( A1 => n1863, A2 => n1296, B1 => n1895, B2 => 
                           n1197, ZN => n4492);
   U2993 : OAI222_X1 port map( A1 => n2151_port, A2 => n1176, B1 => n2183, B2 
                           => n1173, C1 => n2119, C2 => n1170, ZN => n4489);
   U2994 : OAI222_X1 port map( A1 => n2055, A2 => n1185, B1 => n2087, B2 => 
                           n1182, C1 => n2023, C2 => n1179, ZN => n4490);
   U2995 : NOR4_X1 port map( A1 => n4498, A2 => n4499, A3 => n4500, A4 => n4501
                           , ZN => n4497);
   U2996 : OAI22_X1 port map( A1 => n2215, A2 => n782, B1 => n2247, B2 => n779,
                           ZN => n4501);
   U2997 : OAI222_X1 port map( A1 => n2503, A2 => n758, B1 => n2535, B2 => n755
                           , C1 => n2471, C2 => n752, ZN => n4498);
   U2998 : OAI222_X1 port map( A1 => n2407, A2 => n767, B1 => n2439, B2 => n764
                           , C1 => n2375, C2 => n761, ZN => n4499);
   U2999 : NOR4_X1 port map( A1 => n5891, A2 => n5892, A3 => n5893, A4 => n5894
                           , ZN => n5890);
   U3000 : OAI22_X1 port map( A1 => n1862, A2 => n488, B1 => n1894, B2 => n485,
                           ZN => n5894);
   U3001 : OAI222_X1 port map( A1 => n2150, A2 => n464, B1 => n2182, B2 => n461
                           , C1 => n2118, C2 => n458, ZN => n5891);
   U3002 : OAI222_X1 port map( A1 => n2054, A2 => n473, B1 => n2086, B2 => n470
                           , C1 => n2022, C2 => n467, ZN => n5892);
   U3003 : NOR4_X1 port map( A1 => n5900, A2 => n5901, A3 => n5902, A4 => n5903
                           , ZN => n5899);
   U3004 : OAI22_X1 port map( A1 => n2214, A2 => n70, B1 => n2246, B2 => n67, 
                           ZN => n5903);
   U3005 : OAI222_X1 port map( A1 => n2502, A2 => n46, B1 => n2534, B2 => n43, 
                           C1 => n2470, C2 => n40, ZN => n5900);
   U3006 : OAI222_X1 port map( A1 => n2406, A2 => n55, B1 => n2438, B2 => n52, 
                           C1 => n2374, C2 => n49, ZN => n5901);
   U3007 : NOR4_X1 port map( A1 => n4448, A2 => n4449, A3 => n4450, A4 => n4451
                           , ZN => n4447);
   U3008 : OAI22_X1 port map( A1 => n1862, A2 => n1296, B1 => n1894, B2 => 
                           n1197, ZN => n4451);
   U3009 : OAI222_X1 port map( A1 => n2150, A2 => n1176, B1 => n2182, B2 => 
                           n1173, C1 => n2118, C2 => n1170, ZN => n4448);
   U3010 : OAI222_X1 port map( A1 => n2054, A2 => n1185, B1 => n2086, B2 => 
                           n1182, C1 => n2022, C2 => n1179, ZN => n4449);
   U3011 : NOR4_X1 port map( A1 => n4457, A2 => n4458, A3 => n4459, A4 => n4460
                           , ZN => n4456);
   U3012 : OAI22_X1 port map( A1 => n2214, A2 => n782, B1 => n2246, B2 => n779,
                           ZN => n4460);
   U3013 : OAI222_X1 port map( A1 => n2502, A2 => n758, B1 => n2534, B2 => n755
                           , C1 => n2470, C2 => n752, ZN => n4457);
   U3014 : OAI222_X1 port map( A1 => n2406, A2 => n767, B1 => n2438, B2 => n764
                           , C1 => n2374, C2 => n761, ZN => n4458);
   U3015 : NOR4_X1 port map( A1 => n5850, A2 => n5851, A3 => n5852, A4 => n5853
                           , ZN => n5849);
   U3016 : OAI22_X1 port map( A1 => n1861, A2 => n488, B1 => n1893, B2 => n485,
                           ZN => n5853);
   U3017 : OAI222_X1 port map( A1 => n2149, A2 => n464, B1 => n2181, B2 => n461
                           , C1 => n2117, C2 => n458, ZN => n5850);
   U3018 : OAI222_X1 port map( A1 => n2053, A2 => n473, B1 => n2085, B2 => n470
                           , C1 => n2021, C2 => n467, ZN => n5851);
   U3019 : NOR4_X1 port map( A1 => n5859, A2 => n5860, A3 => n5861, A4 => n5862
                           , ZN => n5858);
   U3020 : OAI22_X1 port map( A1 => n2213, A2 => n70, B1 => n2245, B2 => n67, 
                           ZN => n5862);
   U3021 : OAI222_X1 port map( A1 => n2501, A2 => n46, B1 => n2533, B2 => n43, 
                           C1 => n2469, C2 => n40, ZN => n5859);
   U3022 : OAI222_X1 port map( A1 => n2405, A2 => n55, B1 => n2437, B2 => n52, 
                           C1 => n2373, C2 => n49, ZN => n5860);
   U3023 : NOR4_X1 port map( A1 => n4407, A2 => n4408, A3 => n4409, A4 => n4410
                           , ZN => n4406);
   U3024 : OAI22_X1 port map( A1 => n1861, A2 => n1296, B1 => n1893, B2 => 
                           n1197, ZN => n4410);
   U3025 : OAI222_X1 port map( A1 => n2149, A2 => n1176, B1 => n2181, B2 => 
                           n1173, C1 => n2117, C2 => n1170, ZN => n4407);
   U3026 : OAI222_X1 port map( A1 => n2053, A2 => n1185, B1 => n2085, B2 => 
                           n1182, C1 => n2021, C2 => n1179, ZN => n4408);
   U3027 : NOR4_X1 port map( A1 => n4416, A2 => n4417, A3 => n4418, A4 => n4419
                           , ZN => n4415);
   U3028 : OAI22_X1 port map( A1 => n2213, A2 => n782, B1 => n2245, B2 => n779,
                           ZN => n4419);
   U3029 : OAI222_X1 port map( A1 => n2501, A2 => n758, B1 => n2533, B2 => n755
                           , C1 => n2469, C2 => n752, ZN => n4416);
   U3030 : OAI222_X1 port map( A1 => n2405, A2 => n767, B1 => n2437, B2 => n764
                           , C1 => n2373, C2 => n761, ZN => n4417);
   U3031 : NOR4_X1 port map( A1 => n5809, A2 => n5810, A3 => n5811, A4 => n5812
                           , ZN => n5808);
   U3032 : OAI22_X1 port map( A1 => n1860, A2 => n488, B1 => n1892, B2 => n485,
                           ZN => n5812);
   U3033 : OAI222_X1 port map( A1 => n2148, A2 => n464, B1 => n2180, B2 => n461
                           , C1 => n2116, C2 => n458, ZN => n5809);
   U3034 : OAI222_X1 port map( A1 => n2052, A2 => n473, B1 => n2084, B2 => n470
                           , C1 => n2020, C2 => n467, ZN => n5810);
   U3035 : NOR4_X1 port map( A1 => n5818, A2 => n5819, A3 => n5820, A4 => n5821
                           , ZN => n5817);
   U3036 : OAI22_X1 port map( A1 => n2212, A2 => n70, B1 => n2244, B2 => n67, 
                           ZN => n5821);
   U3037 : OAI222_X1 port map( A1 => n2500, A2 => n46, B1 => n2532, B2 => n43, 
                           C1 => n2468, C2 => n40, ZN => n5818);
   U3038 : OAI222_X1 port map( A1 => n2404, A2 => n55, B1 => n2436, B2 => n52, 
                           C1 => n2372, C2 => n49, ZN => n5819);
   U3039 : NOR4_X1 port map( A1 => n4366, A2 => n4367, A3 => n4368, A4 => n4369
                           , ZN => n4365);
   U3040 : OAI22_X1 port map( A1 => n1860, A2 => n1296, B1 => n1892, B2 => 
                           n1197, ZN => n4369);
   U3041 : OAI222_X1 port map( A1 => n2148, A2 => n1176, B1 => n2180, B2 => 
                           n1173, C1 => n2116, C2 => n1170, ZN => n4366);
   U3042 : OAI222_X1 port map( A1 => n2052, A2 => n1185, B1 => n2084, B2 => 
                           n1182, C1 => n2020, C2 => n1179, ZN => n4367);
   U3043 : NOR4_X1 port map( A1 => n4375, A2 => n4376, A3 => n4377, A4 => n4378
                           , ZN => n4374);
   U3044 : OAI22_X1 port map( A1 => n2212, A2 => n782, B1 => n2244, B2 => n779,
                           ZN => n4378);
   U3045 : OAI222_X1 port map( A1 => n2500, A2 => n758, B1 => n2532, B2 => n755
                           , C1 => n2468, C2 => n752, ZN => n4375);
   U3046 : OAI222_X1 port map( A1 => n2404, A2 => n767, B1 => n2436, B2 => n764
                           , C1 => n2372, C2 => n761, ZN => n4376);
   U3047 : NOR4_X1 port map( A1 => n5768, A2 => n5769, A3 => n5770, A4 => n5771
                           , ZN => n5767);
   U3048 : OAI22_X1 port map( A1 => n1859, A2 => n489, B1 => n1891, B2 => n486,
                           ZN => n5771);
   U3049 : OAI222_X1 port map( A1 => n2147, A2 => n465, B1 => n2179, B2 => n462
                           , C1 => n2115, C2 => n459, ZN => n5768);
   U3050 : OAI222_X1 port map( A1 => n2051, A2 => n474, B1 => n2083, B2 => n471
                           , C1 => n2019, C2 => n468, ZN => n5769);
   U3051 : NOR4_X1 port map( A1 => n5777, A2 => n5778, A3 => n5779, A4 => n5780
                           , ZN => n5776);
   U3052 : OAI22_X1 port map( A1 => n2211, A2 => n71, B1 => n2243, B2 => n68, 
                           ZN => n5780);
   U3053 : OAI222_X1 port map( A1 => n2499, A2 => n47, B1 => n2531, B2 => n44, 
                           C1 => n2467, C2 => n41, ZN => n5777);
   U3054 : OAI222_X1 port map( A1 => n2403, A2 => n56, B1 => n2435, B2 => n53, 
                           C1 => n2371, C2 => n50, ZN => n5778);
   U3055 : NOR4_X1 port map( A1 => n4325, A2 => n4326, A3 => n4327, A4 => n4328
                           , ZN => n4324);
   U3056 : OAI22_X1 port map( A1 => n1859, A2 => n1297, B1 => n1891, B2 => 
                           n1198, ZN => n4328);
   U3057 : OAI222_X1 port map( A1 => n2147, A2 => n1177, B1 => n2179, B2 => 
                           n1174, C1 => n2115, C2 => n1171, ZN => n4325);
   U3058 : OAI222_X1 port map( A1 => n2051, A2 => n1186, B1 => n2083, B2 => 
                           n1183, C1 => n2019, C2 => n1180, ZN => n4326);
   U3059 : NOR4_X1 port map( A1 => n4334, A2 => n4335, A3 => n4336, A4 => n4337
                           , ZN => n4333);
   U3060 : OAI22_X1 port map( A1 => n2211, A2 => n783, B1 => n2243, B2 => n780,
                           ZN => n4337);
   U3061 : OAI222_X1 port map( A1 => n2499, A2 => n759, B1 => n2531, B2 => n756
                           , C1 => n2467, C2 => n753, ZN => n4334);
   U3062 : OAI222_X1 port map( A1 => n2403, A2 => n768, B1 => n2435, B2 => n765
                           , C1 => n2371, C2 => n762, ZN => n4335);
   U3063 : NOR4_X1 port map( A1 => n5727, A2 => n5728, A3 => n5729, A4 => n5730
                           , ZN => n5726);
   U3064 : OAI22_X1 port map( A1 => n1858, A2 => n489, B1 => n1890, B2 => n486,
                           ZN => n5730);
   U3065 : OAI222_X1 port map( A1 => n2146, A2 => n465, B1 => n2178, B2 => n462
                           , C1 => n2114, C2 => n459, ZN => n5727);
   U3066 : OAI222_X1 port map( A1 => n2050, A2 => n474, B1 => n2082, B2 => n471
                           , C1 => n2018, C2 => n468, ZN => n5728);
   U3067 : NOR4_X1 port map( A1 => n5736, A2 => n5737, A3 => n5738, A4 => n5739
                           , ZN => n5735);
   U3068 : OAI22_X1 port map( A1 => n2210, A2 => n71, B1 => n2242, B2 => n68, 
                           ZN => n5739);
   U3069 : OAI222_X1 port map( A1 => n2498, A2 => n47, B1 => n2530, B2 => n44, 
                           C1 => n2466, C2 => n41, ZN => n5736);
   U3070 : OAI222_X1 port map( A1 => n2402, A2 => n56, B1 => n2434, B2 => n53, 
                           C1 => n2370, C2 => n50, ZN => n5737);
   U3071 : NOR4_X1 port map( A1 => n4284, A2 => n4285, A3 => n4286, A4 => n4287
                           , ZN => n4283);
   U3072 : OAI22_X1 port map( A1 => n1858, A2 => n1297, B1 => n1890, B2 => 
                           n1198, ZN => n4287);
   U3073 : OAI222_X1 port map( A1 => n2146, A2 => n1177, B1 => n2178, B2 => 
                           n1174, C1 => n2114, C2 => n1171, ZN => n4284);
   U3074 : OAI222_X1 port map( A1 => n2050, A2 => n1186, B1 => n2082, B2 => 
                           n1183, C1 => n2018, C2 => n1180, ZN => n4285);
   U3075 : NOR4_X1 port map( A1 => n4293, A2 => n4294, A3 => n4295, A4 => n4296
                           , ZN => n4292);
   U3076 : OAI22_X1 port map( A1 => n2210, A2 => n783, B1 => n2242, B2 => n780,
                           ZN => n4296);
   U3077 : OAI222_X1 port map( A1 => n2498, A2 => n759, B1 => n2530, B2 => n756
                           , C1 => n2466, C2 => n753, ZN => n4293);
   U3078 : OAI222_X1 port map( A1 => n2402, A2 => n768, B1 => n2434, B2 => n765
                           , C1 => n2370, C2 => n762, ZN => n4294);
   U3079 : NOR4_X1 port map( A1 => n5686, A2 => n5687, A3 => n5688, A4 => n5689
                           , ZN => n5685);
   U3080 : OAI22_X1 port map( A1 => n1857, A2 => n489, B1 => n1889, B2 => n486,
                           ZN => n5689);
   U3081 : OAI222_X1 port map( A1 => n2145, A2 => n465, B1 => n2177, B2 => n462
                           , C1 => n2113, C2 => n459, ZN => n5686);
   U3082 : OAI222_X1 port map( A1 => n2049, A2 => n474, B1 => n2081, B2 => n471
                           , C1 => n2017, C2 => n468, ZN => n5687);
   U3083 : NOR4_X1 port map( A1 => n5695, A2 => n5696, A3 => n5697, A4 => n5698
                           , ZN => n5694);
   U3084 : OAI22_X1 port map( A1 => n2209, A2 => n71, B1 => n2241, B2 => n68, 
                           ZN => n5698);
   U3085 : OAI222_X1 port map( A1 => n2497, A2 => n47, B1 => n2529, B2 => n44, 
                           C1 => n2465, C2 => n41, ZN => n5695);
   U3086 : OAI222_X1 port map( A1 => n2401, A2 => n56, B1 => n2433, B2 => n53, 
                           C1 => n2369, C2 => n50, ZN => n5696);
   U3087 : NOR4_X1 port map( A1 => n4243, A2 => n4244, A3 => n4245, A4 => n4246
                           , ZN => n4242);
   U3088 : OAI22_X1 port map( A1 => n1857, A2 => n1297, B1 => n1889, B2 => 
                           n1198, ZN => n4246);
   U3089 : OAI222_X1 port map( A1 => n2145, A2 => n1177, B1 => n2177, B2 => 
                           n1174, C1 => n2113, C2 => n1171, ZN => n4243);
   U3090 : OAI222_X1 port map( A1 => n2049, A2 => n1186, B1 => n2081, B2 => 
                           n1183, C1 => n2017, C2 => n1180, ZN => n4244);
   U3091 : NOR4_X1 port map( A1 => n4252, A2 => n4253, A3 => n4254, A4 => n4255
                           , ZN => n4251);
   U3092 : OAI22_X1 port map( A1 => n2209, A2 => n783, B1 => n2241, B2 => n780,
                           ZN => n4255);
   U3093 : OAI222_X1 port map( A1 => n2497, A2 => n759, B1 => n2529, B2 => n756
                           , C1 => n2465, C2 => n753, ZN => n4252);
   U3094 : OAI222_X1 port map( A1 => n2401, A2 => n768, B1 => n2433, B2 => n765
                           , C1 => n2369, C2 => n762, ZN => n4253);
   U3095 : NOR4_X1 port map( A1 => n5645, A2 => n5646, A3 => n5647, A4 => n5648
                           , ZN => n5644);
   U3096 : OAI22_X1 port map( A1 => n1856, A2 => n489, B1 => n1888, B2 => n486,
                           ZN => n5648);
   U3097 : OAI222_X1 port map( A1 => n2144, A2 => n465, B1 => n2176, B2 => n462
                           , C1 => n2112, C2 => n459, ZN => n5645);
   U3098 : OAI222_X1 port map( A1 => n2048, A2 => n474, B1 => n2080, B2 => n471
                           , C1 => n2016, C2 => n468, ZN => n5646);
   U3099 : NOR4_X1 port map( A1 => n5654, A2 => n5655, A3 => n5656, A4 => n5657
                           , ZN => n5653);
   U3100 : OAI22_X1 port map( A1 => n2208, A2 => n71, B1 => n2240, B2 => n68, 
                           ZN => n5657);
   U3101 : OAI222_X1 port map( A1 => n2496, A2 => n47, B1 => n2528, B2 => n44, 
                           C1 => n2464, C2 => n41, ZN => n5654);
   U3102 : OAI222_X1 port map( A1 => n2400, A2 => n56, B1 => n2432, B2 => n53, 
                           C1 => n2368, C2 => n50, ZN => n5655);
   U3103 : NOR4_X1 port map( A1 => n4202, A2 => n4203, A3 => n4204, A4 => n4205
                           , ZN => n4201);
   U3104 : OAI22_X1 port map( A1 => n1856, A2 => n1297, B1 => n1888, B2 => 
                           n1198, ZN => n4205);
   U3105 : OAI222_X1 port map( A1 => n2144, A2 => n1177, B1 => n2176, B2 => 
                           n1174, C1 => n2112, C2 => n1171, ZN => n4202);
   U3106 : OAI222_X1 port map( A1 => n2048, A2 => n1186, B1 => n2080, B2 => 
                           n1183, C1 => n2016, C2 => n1180, ZN => n4203);
   U3107 : NOR4_X1 port map( A1 => n4211, A2 => n4212, A3 => n4213, A4 => n4214
                           , ZN => n4210);
   U3108 : OAI22_X1 port map( A1 => n2208, A2 => n783, B1 => n2240, B2 => n780,
                           ZN => n4214);
   U3109 : OAI222_X1 port map( A1 => n2496, A2 => n759, B1 => n2528, B2 => n756
                           , C1 => n2464, C2 => n753, ZN => n4211);
   U3110 : OAI222_X1 port map( A1 => n2400, A2 => n768, B1 => n2432, B2 => n765
                           , C1 => n2368, C2 => n762, ZN => n4212);
   U3111 : NOR4_X1 port map( A1 => n5604, A2 => n5605, A3 => n5606, A4 => n5607
                           , ZN => n5603);
   U3112 : OAI22_X1 port map( A1 => n1855, A2 => n489, B1 => n1887, B2 => n486,
                           ZN => n5607);
   U3113 : OAI222_X1 port map( A1 => n2143, A2 => n465, B1 => n2175, B2 => n462
                           , C1 => n2111, C2 => n459, ZN => n5604);
   U3114 : OAI222_X1 port map( A1 => n2047, A2 => n474, B1 => n2079, B2 => n471
                           , C1 => n2015, C2 => n468, ZN => n5605);
   U3115 : NOR4_X1 port map( A1 => n5613, A2 => n5614, A3 => n5615, A4 => n5616
                           , ZN => n5612);
   U3116 : OAI22_X1 port map( A1 => n2207, A2 => n71, B1 => n2239, B2 => n68, 
                           ZN => n5616);
   U3117 : OAI222_X1 port map( A1 => n2495, A2 => n47, B1 => n2527, B2 => n44, 
                           C1 => n2463, C2 => n41, ZN => n5613);
   U3118 : OAI222_X1 port map( A1 => n2399, A2 => n56, B1 => n2431, B2 => n53, 
                           C1 => n2367, C2 => n50, ZN => n5614);
   U3119 : NOR4_X1 port map( A1 => n4161, A2 => n4162, A3 => n4163, A4 => n4164
                           , ZN => n4160);
   U3120 : OAI22_X1 port map( A1 => n1855, A2 => n1297, B1 => n1887, B2 => 
                           n1198, ZN => n4164);
   U3121 : OAI222_X1 port map( A1 => n2143, A2 => n1177, B1 => n2175, B2 => 
                           n1174, C1 => n2111, C2 => n1171, ZN => n4161);
   U3122 : OAI222_X1 port map( A1 => n2047, A2 => n1186, B1 => n2079, B2 => 
                           n1183, C1 => n2015, C2 => n1180, ZN => n4162);
   U3123 : NOR4_X1 port map( A1 => n4170, A2 => n4171, A3 => n4172, A4 => n4173
                           , ZN => n4169);
   U3124 : OAI22_X1 port map( A1 => n2207, A2 => n783, B1 => n2239, B2 => n780,
                           ZN => n4173);
   U3125 : OAI222_X1 port map( A1 => n2495, A2 => n759, B1 => n2527, B2 => n756
                           , C1 => n2463, C2 => n753, ZN => n4170);
   U3126 : OAI222_X1 port map( A1 => n2399, A2 => n768, B1 => n2431, B2 => n765
                           , C1 => n2367, C2 => n762, ZN => n4171);
   U3127 : NOR4_X1 port map( A1 => n5563, A2 => n5564, A3 => n5565, A4 => n5566
                           , ZN => n5562);
   U3128 : OAI22_X1 port map( A1 => n1854, A2 => n489, B1 => n1886, B2 => n486,
                           ZN => n5566);
   U3129 : OAI222_X1 port map( A1 => n2142, A2 => n465, B1 => n2174, B2 => n462
                           , C1 => n2110, C2 => n459, ZN => n5563);
   U3130 : OAI222_X1 port map( A1 => n2046, A2 => n474, B1 => n2078, B2 => n471
                           , C1 => n2014, C2 => n468, ZN => n5564);
   U3131 : NOR4_X1 port map( A1 => n5572, A2 => n5573, A3 => n5574, A4 => n5575
                           , ZN => n5571);
   U3132 : OAI22_X1 port map( A1 => n2206, A2 => n71, B1 => n2238, B2 => n68, 
                           ZN => n5575);
   U3133 : OAI222_X1 port map( A1 => n2494, A2 => n47, B1 => n2526, B2 => n44, 
                           C1 => n2462, C2 => n41, ZN => n5572);
   U3134 : OAI222_X1 port map( A1 => n2398, A2 => n56, B1 => n2430, B2 => n53, 
                           C1 => n2366, C2 => n50, ZN => n5573);
   U3135 : NOR4_X1 port map( A1 => n4120, A2 => n4121, A3 => n4122, A4 => n4123
                           , ZN => n4119);
   U3136 : OAI22_X1 port map( A1 => n1854, A2 => n1297, B1 => n1886, B2 => 
                           n1198, ZN => n4123);
   U3137 : OAI222_X1 port map( A1 => n2142, A2 => n1177, B1 => n2174, B2 => 
                           n1174, C1 => n2110, C2 => n1171, ZN => n4120);
   U3138 : OAI222_X1 port map( A1 => n2046, A2 => n1186, B1 => n2078, B2 => 
                           n1183, C1 => n2014, C2 => n1180, ZN => n4121);
   U3139 : NOR4_X1 port map( A1 => n4129, A2 => n4130, A3 => n4131, A4 => n4132
                           , ZN => n4128);
   U3140 : OAI22_X1 port map( A1 => n2206, A2 => n783, B1 => n2238, B2 => n780,
                           ZN => n4132);
   U3141 : OAI222_X1 port map( A1 => n2494, A2 => n759, B1 => n2526, B2 => n756
                           , C1 => n2462, C2 => n753, ZN => n4129);
   U3142 : OAI222_X1 port map( A1 => n2398, A2 => n768, B1 => n2430, B2 => n765
                           , C1 => n2366, C2 => n762, ZN => n4130);
   U3143 : NOR4_X1 port map( A1 => n5522, A2 => n5523, A3 => n5524, A4 => n5525
                           , ZN => n5521);
   U3144 : OAI22_X1 port map( A1 => n1853, A2 => n489, B1 => n1885, B2 => n486,
                           ZN => n5525);
   U3145 : OAI222_X1 port map( A1 => n2141, A2 => n465, B1 => n2173, B2 => n462
                           , C1 => n2109, C2 => n459, ZN => n5522);
   U3146 : OAI222_X1 port map( A1 => n2045, A2 => n474, B1 => n2077, B2 => n471
                           , C1 => n2013, C2 => n468, ZN => n5523);
   U3147 : NOR4_X1 port map( A1 => n5531, A2 => n5532, A3 => n5533, A4 => n5534
                           , ZN => n5530);
   U3148 : OAI22_X1 port map( A1 => n2205, A2 => n71, B1 => n2237, B2 => n68, 
                           ZN => n5534);
   U3149 : OAI222_X1 port map( A1 => n2493, A2 => n47, B1 => n2525, B2 => n44, 
                           C1 => n2461, C2 => n41, ZN => n5531);
   U3150 : OAI222_X1 port map( A1 => n2397, A2 => n56, B1 => n2429, B2 => n53, 
                           C1 => n2365, C2 => n50, ZN => n5532);
   U3151 : NOR4_X1 port map( A1 => n4079, A2 => n4080, A3 => n4081, A4 => n4082
                           , ZN => n4078);
   U3152 : OAI22_X1 port map( A1 => n1853, A2 => n1297, B1 => n1885, B2 => 
                           n1198, ZN => n4082);
   U3153 : OAI222_X1 port map( A1 => n2141, A2 => n1177, B1 => n2173, B2 => 
                           n1174, C1 => n2109, C2 => n1171, ZN => n4079);
   U3154 : OAI222_X1 port map( A1 => n2045, A2 => n1186, B1 => n2077, B2 => 
                           n1183, C1 => n2013, C2 => n1180, ZN => n4080);
   U3155 : NOR4_X1 port map( A1 => n4088, A2 => n4089, A3 => n4090, A4 => n4091
                           , ZN => n4087);
   U3156 : OAI22_X1 port map( A1 => n2205, A2 => n783, B1 => n2237, B2 => n780,
                           ZN => n4091);
   U3157 : OAI222_X1 port map( A1 => n2493, A2 => n759, B1 => n2525, B2 => n756
                           , C1 => n2461, C2 => n753, ZN => n4088);
   U3158 : OAI222_X1 port map( A1 => n2397, A2 => n768, B1 => n2429, B2 => n765
                           , C1 => n2365, C2 => n762, ZN => n4089);
   U3159 : NOR4_X1 port map( A1 => n5481, A2 => n5482, A3 => n5483, A4 => n5484
                           , ZN => n5480);
   U3160 : OAI22_X1 port map( A1 => n1852, A2 => n489, B1 => n1884, B2 => n486,
                           ZN => n5484);
   U3161 : OAI222_X1 port map( A1 => n2140, A2 => n465, B1 => n2172, B2 => n462
                           , C1 => n2108, C2 => n459, ZN => n5481);
   U3162 : OAI222_X1 port map( A1 => n2044, A2 => n474, B1 => n2076, B2 => n471
                           , C1 => n2012, C2 => n468, ZN => n5482);
   U3163 : NOR4_X1 port map( A1 => n5490, A2 => n5491, A3 => n5492, A4 => n5493
                           , ZN => n5489);
   U3164 : OAI22_X1 port map( A1 => n2204, A2 => n71, B1 => n2236, B2 => n68, 
                           ZN => n5493);
   U3165 : OAI222_X1 port map( A1 => n2492, A2 => n47, B1 => n2524, B2 => n44, 
                           C1 => n2460, C2 => n41, ZN => n5490);
   U3166 : OAI222_X1 port map( A1 => n2396, A2 => n56, B1 => n2428, B2 => n53, 
                           C1 => n2364, C2 => n50, ZN => n5491);
   U3167 : NOR4_X1 port map( A1 => n4038, A2 => n4039, A3 => n4040, A4 => n4041
                           , ZN => n4037);
   U3168 : OAI22_X1 port map( A1 => n1852, A2 => n1297, B1 => n1884, B2 => 
                           n1198, ZN => n4041);
   U3169 : OAI222_X1 port map( A1 => n2140, A2 => n1177, B1 => n2172, B2 => 
                           n1174, C1 => n2108, C2 => n1171, ZN => n4038);
   U3170 : OAI222_X1 port map( A1 => n2044, A2 => n1186, B1 => n2076, B2 => 
                           n1183, C1 => n2012, C2 => n1180, ZN => n4039);
   U3171 : NOR4_X1 port map( A1 => n4047, A2 => n4048, A3 => n4049, A4 => n4050
                           , ZN => n4046);
   U3172 : OAI22_X1 port map( A1 => n2204, A2 => n783, B1 => n2236, B2 => n780,
                           ZN => n4050);
   U3173 : OAI222_X1 port map( A1 => n2492, A2 => n759, B1 => n2524, B2 => n756
                           , C1 => n2460, C2 => n753, ZN => n4047);
   U3174 : OAI222_X1 port map( A1 => n2396, A2 => n768, B1 => n2428, B2 => n765
                           , C1 => n2364, C2 => n762, ZN => n4048);
   U3175 : NOR4_X1 port map( A1 => n5440, A2 => n5441, A3 => n5442, A4 => n5443
                           , ZN => n5439);
   U3176 : OAI22_X1 port map( A1 => n1851, A2 => n489, B1 => n1883, B2 => n486,
                           ZN => n5443);
   U3177 : OAI222_X1 port map( A1 => n2139, A2 => n465, B1 => n2171, B2 => n462
                           , C1 => n2107, C2 => n459, ZN => n5440);
   U3178 : OAI222_X1 port map( A1 => n2043, A2 => n474, B1 => n2075, B2 => n471
                           , C1 => n2011, C2 => n468, ZN => n5441);
   U3179 : NOR4_X1 port map( A1 => n5449, A2 => n5450, A3 => n5451, A4 => n5452
                           , ZN => n5448);
   U3180 : OAI22_X1 port map( A1 => n2203, A2 => n71, B1 => n2235, B2 => n68, 
                           ZN => n5452);
   U3181 : OAI222_X1 port map( A1 => n2491, A2 => n47, B1 => n2523, B2 => n44, 
                           C1 => n2459, C2 => n41, ZN => n5449);
   U3182 : OAI222_X1 port map( A1 => n2395, A2 => n56, B1 => n2427, B2 => n53, 
                           C1 => n2363, C2 => n50, ZN => n5450);
   U3183 : NOR4_X1 port map( A1 => n3997, A2 => n3998, A3 => n3999, A4 => n4000
                           , ZN => n3996);
   U3184 : OAI22_X1 port map( A1 => n1851, A2 => n1297, B1 => n1883, B2 => 
                           n1198, ZN => n4000);
   U3185 : OAI222_X1 port map( A1 => n2139, A2 => n1177, B1 => n2171, B2 => 
                           n1174, C1 => n2107, C2 => n1171, ZN => n3997);
   U3186 : OAI222_X1 port map( A1 => n2043, A2 => n1186, B1 => n2075, B2 => 
                           n1183, C1 => n2011, C2 => n1180, ZN => n3998);
   U3187 : NOR4_X1 port map( A1 => n4006, A2 => n4007, A3 => n4008, A4 => n4009
                           , ZN => n4005);
   U3188 : OAI22_X1 port map( A1 => n2203, A2 => n783, B1 => n2235, B2 => n780,
                           ZN => n4009);
   U3189 : OAI222_X1 port map( A1 => n2491, A2 => n759, B1 => n2523, B2 => n756
                           , C1 => n2459, C2 => n753, ZN => n4006);
   U3190 : OAI222_X1 port map( A1 => n2395, A2 => n768, B1 => n2427, B2 => n765
                           , C1 => n2363, C2 => n762, ZN => n4007);
   U3191 : NOR4_X1 port map( A1 => n5399, A2 => n5400, A3 => n5401, A4 => n5402
                           , ZN => n5398);
   U3192 : OAI22_X1 port map( A1 => n1850, A2 => n489, B1 => n1882, B2 => n486,
                           ZN => n5402);
   U3193 : OAI222_X1 port map( A1 => n2138, A2 => n465, B1 => n2170, B2 => n462
                           , C1 => n2106, C2 => n459, ZN => n5399);
   U3194 : OAI222_X1 port map( A1 => n2042, A2 => n474, B1 => n2074, B2 => n471
                           , C1 => n2010, C2 => n468, ZN => n5400);
   U3195 : NOR4_X1 port map( A1 => n5408, A2 => n5409, A3 => n5410, A4 => n5411
                           , ZN => n5407);
   U3196 : OAI22_X1 port map( A1 => n2202, A2 => n71, B1 => n2234, B2 => n68, 
                           ZN => n5411);
   U3197 : OAI222_X1 port map( A1 => n2490, A2 => n47, B1 => n2522, B2 => n44, 
                           C1 => n2458, C2 => n41, ZN => n5408);
   U3198 : OAI222_X1 port map( A1 => n2394, A2 => n56, B1 => n2426, B2 => n53, 
                           C1 => n2362, C2 => n50, ZN => n5409);
   U3199 : NOR4_X1 port map( A1 => n3956, A2 => n3957, A3 => n3958, A4 => n3959
                           , ZN => n3955);
   U3200 : OAI22_X1 port map( A1 => n1850, A2 => n1297, B1 => n1882, B2 => 
                           n1198, ZN => n3959);
   U3201 : OAI222_X1 port map( A1 => n2138, A2 => n1177, B1 => n2170, B2 => 
                           n1174, C1 => n2106, C2 => n1171, ZN => n3956);
   U3202 : OAI222_X1 port map( A1 => n2042, A2 => n1186, B1 => n2074, B2 => 
                           n1183, C1 => n2010, C2 => n1180, ZN => n3957);
   U3203 : NOR4_X1 port map( A1 => n3965, A2 => n3966, A3 => n3967, A4 => n3968
                           , ZN => n3964);
   U3204 : OAI22_X1 port map( A1 => n2202, A2 => n783, B1 => n2234, B2 => n780,
                           ZN => n3968);
   U3205 : OAI222_X1 port map( A1 => n2490, A2 => n759, B1 => n2522, B2 => n756
                           , C1 => n2458, C2 => n753, ZN => n3965);
   U3206 : OAI222_X1 port map( A1 => n2394, A2 => n768, B1 => n2426, B2 => n765
                           , C1 => n2362, C2 => n762, ZN => n3966);
   U3207 : NOR4_X1 port map( A1 => n5358, A2 => n5359, A3 => n5360, A4 => n5361
                           , ZN => n5357);
   U3208 : OAI22_X1 port map( A1 => n1849, A2 => n489, B1 => n1881, B2 => n486,
                           ZN => n5361);
   U3209 : OAI222_X1 port map( A1 => n2137, A2 => n465, B1 => n2169, B2 => n462
                           , C1 => n2105, C2 => n459, ZN => n5358);
   U3210 : OAI222_X1 port map( A1 => n2041, A2 => n474, B1 => n2073, B2 => n471
                           , C1 => n2009, C2 => n468, ZN => n5359);
   U3211 : NOR4_X1 port map( A1 => n5367, A2 => n5368, A3 => n5369, A4 => n5370
                           , ZN => n5366);
   U3212 : OAI22_X1 port map( A1 => n2201, A2 => n71, B1 => n2233, B2 => n68, 
                           ZN => n5370);
   U3213 : OAI222_X1 port map( A1 => n2489, A2 => n47, B1 => n2521, B2 => n44, 
                           C1 => n2457, C2 => n41, ZN => n5367);
   U3214 : OAI222_X1 port map( A1 => n2393, A2 => n56, B1 => n2425, B2 => n53, 
                           C1 => n2361, C2 => n50, ZN => n5368);
   U3215 : NOR4_X1 port map( A1 => n3915, A2 => n3916, A3 => n3917, A4 => n3918
                           , ZN => n3914);
   U3216 : OAI22_X1 port map( A1 => n1849, A2 => n1297, B1 => n1881, B2 => 
                           n1198, ZN => n3918);
   U3217 : OAI222_X1 port map( A1 => n2137, A2 => n1177, B1 => n2169, B2 => 
                           n1174, C1 => n2105, C2 => n1171, ZN => n3915);
   U3218 : OAI222_X1 port map( A1 => n2041, A2 => n1186, B1 => n2073, B2 => 
                           n1183, C1 => n2009, C2 => n1180, ZN => n3916);
   U3219 : NOR4_X1 port map( A1 => n3924, A2 => n3925, A3 => n3926, A4 => n3927
                           , ZN => n3923);
   U3220 : OAI22_X1 port map( A1 => n2201, A2 => n783, B1 => n2233, B2 => n780,
                           ZN => n3927);
   U3221 : OAI222_X1 port map( A1 => n2489, A2 => n759, B1 => n2521, B2 => n756
                           , C1 => n2457, C2 => n753, ZN => n3924);
   U3222 : OAI222_X1 port map( A1 => n2393, A2 => n768, B1 => n2425, B2 => n765
                           , C1 => n2361, C2 => n762, ZN => n3925);
   U3223 : NOR4_X1 port map( A1 => n5317, A2 => n5318, A3 => n5319, A4 => n5320
                           , ZN => n5316);
   U3224 : OAI22_X1 port map( A1 => n1848, A2 => n489, B1 => n1880, B2 => n486,
                           ZN => n5320);
   U3225 : OAI222_X1 port map( A1 => n2136, A2 => n465, B1 => n2168, B2 => n462
                           , C1 => n2104, C2 => n459, ZN => n5317);
   U3226 : OAI222_X1 port map( A1 => n2040, A2 => n474, B1 => n2072, B2 => n471
                           , C1 => n2008, C2 => n468, ZN => n5318);
   U3227 : NOR4_X1 port map( A1 => n5326, A2 => n5327, A3 => n5328, A4 => n5329
                           , ZN => n5325);
   U3228 : OAI22_X1 port map( A1 => n2200, A2 => n71, B1 => n2232, B2 => n68, 
                           ZN => n5329);
   U3229 : OAI222_X1 port map( A1 => n2488, A2 => n47, B1 => n2520, B2 => n44, 
                           C1 => n2456, C2 => n41, ZN => n5326);
   U3230 : OAI222_X1 port map( A1 => n2392, A2 => n56, B1 => n2424, B2 => n53, 
                           C1 => n2360, C2 => n50, ZN => n5327);
   U3231 : NOR4_X1 port map( A1 => n3874, A2 => n3875, A3 => n3876, A4 => n3877
                           , ZN => n3873);
   U3232 : OAI22_X1 port map( A1 => n1848, A2 => n1297, B1 => n1880, B2 => 
                           n1198, ZN => n3877);
   U3233 : OAI222_X1 port map( A1 => n2136, A2 => n1177, B1 => n2168, B2 => 
                           n1174, C1 => n2104, C2 => n1171, ZN => n3874);
   U3234 : OAI222_X1 port map( A1 => n2040, A2 => n1186, B1 => n2072, B2 => 
                           n1183, C1 => n2008, C2 => n1180, ZN => n3875);
   U3235 : NOR4_X1 port map( A1 => n3883, A2 => n3884, A3 => n3885, A4 => n3886
                           , ZN => n3882);
   U3236 : OAI22_X1 port map( A1 => n2200, A2 => n783, B1 => n2232, B2 => n780,
                           ZN => n3886);
   U3237 : OAI222_X1 port map( A1 => n2488, A2 => n759, B1 => n2520, B2 => n756
                           , C1 => n2456, C2 => n753, ZN => n3883);
   U3238 : OAI222_X1 port map( A1 => n2392, A2 => n768, B1 => n2424, B2 => n765
                           , C1 => n2360, C2 => n762, ZN => n3884);
   U3239 : NOR4_X1 port map( A1 => n5276, A2 => n5277, A3 => n5278, A4 => n5279
                           , ZN => n5275);
   U3240 : OAI22_X1 port map( A1 => n1847, A2 => n490, B1 => n1879, B2 => n487,
                           ZN => n5279);
   U3241 : OAI222_X1 port map( A1 => n2135, A2 => n466, B1 => n2167, B2 => n463
                           , C1 => n2103, C2 => n460, ZN => n5276);
   U3242 : OAI222_X1 port map( A1 => n2039, A2 => n475, B1 => n2071, B2 => n472
                           , C1 => n2007, C2 => n469, ZN => n5277);
   U3243 : NOR4_X1 port map( A1 => n5285, A2 => n5286, A3 => n5287, A4 => n5288
                           , ZN => n5284);
   U3244 : OAI22_X1 port map( A1 => n2199, A2 => n72, B1 => n2231, B2 => n69, 
                           ZN => n5288);
   U3245 : OAI222_X1 port map( A1 => n2487, A2 => n48, B1 => n2519, B2 => n45, 
                           C1 => n2455, C2 => n42, ZN => n5285);
   U3246 : OAI222_X1 port map( A1 => n2391, A2 => n57, B1 => n2423, B2 => n54, 
                           C1 => n2359, C2 => n51, ZN => n5286);
   U3247 : NOR4_X1 port map( A1 => n3833, A2 => n3834, A3 => n3835, A4 => n3836
                           , ZN => n3832);
   U3248 : OAI22_X1 port map( A1 => n1847, A2 => n1298, B1 => n1879, B2 => 
                           n1199, ZN => n3836);
   U3249 : OAI222_X1 port map( A1 => n2135, A2 => n1178, B1 => n2167, B2 => 
                           n1175, C1 => n2103, C2 => n1172, ZN => n3833);
   U3250 : OAI222_X1 port map( A1 => n2039, A2 => n1187, B1 => n2071, B2 => 
                           n1184, C1 => n2007, C2 => n1181, ZN => n3834);
   U3251 : NOR4_X1 port map( A1 => n3842, A2 => n3843, A3 => n3844, A4 => n3845
                           , ZN => n3841);
   U3252 : OAI22_X1 port map( A1 => n2199, A2 => n1136, B1 => n2231, B2 => n781
                           , ZN => n3845);
   U3253 : OAI222_X1 port map( A1 => n2487, A2 => n760, B1 => n2519, B2 => n757
                           , C1 => n2455, C2 => n754, ZN => n3842);
   U3254 : OAI222_X1 port map( A1 => n2391, A2 => n769, B1 => n2423, B2 => n766
                           , C1 => n2359, C2 => n763, ZN => n3843);
   U3255 : NOR4_X1 port map( A1 => n5235, A2 => n5236, A3 => n5237, A4 => n5238
                           , ZN => n5234);
   U3256 : OAI22_X1 port map( A1 => n1846, A2 => n490, B1 => n1878, B2 => n487,
                           ZN => n5238);
   U3257 : OAI222_X1 port map( A1 => n2134, A2 => n466, B1 => n2166_port, B2 =>
                           n463, C1 => n2102, C2 => n460, ZN => n5235);
   U3258 : OAI222_X1 port map( A1 => n2038, A2 => n475, B1 => n2070, B2 => n472
                           , C1 => n2006, C2 => n469, ZN => n5236);
   U3259 : NOR4_X1 port map( A1 => n5244, A2 => n5245, A3 => n5246, A4 => n5247
                           , ZN => n5243);
   U3260 : OAI22_X1 port map( A1 => n2198, A2 => n72, B1 => n2230, B2 => n69, 
                           ZN => n5247);
   U3261 : OAI222_X1 port map( A1 => n2486, A2 => n48, B1 => n2518, B2 => n45, 
                           C1 => n2454, C2 => n42, ZN => n5244);
   U3262 : OAI222_X1 port map( A1 => n2390, A2 => n57, B1 => n2422, B2 => n54, 
                           C1 => n2358, C2 => n51, ZN => n5245);
   U3263 : NOR4_X1 port map( A1 => n3792, A2 => n3793, A3 => n3794, A4 => n3795
                           , ZN => n3791);
   U3264 : OAI22_X1 port map( A1 => n1846, A2 => n1298, B1 => n1878, B2 => 
                           n1199, ZN => n3795);
   U3265 : OAI222_X1 port map( A1 => n2134, A2 => n1178, B1 => n2166_port, B2 
                           => n1175, C1 => n2102, C2 => n1172, ZN => n3792);
   U3266 : OAI222_X1 port map( A1 => n2038, A2 => n1187, B1 => n2070, B2 => 
                           n1184, C1 => n2006, C2 => n1181, ZN => n3793);
   U3267 : NOR4_X1 port map( A1 => n3801, A2 => n3802, A3 => n3803, A4 => n3804
                           , ZN => n3800);
   U3268 : OAI22_X1 port map( A1 => n2198, A2 => n1136, B1 => n2230, B2 => n781
                           , ZN => n3804);
   U3269 : OAI222_X1 port map( A1 => n2486, A2 => n760, B1 => n2518, B2 => n757
                           , C1 => n2454, C2 => n754, ZN => n3801);
   U3270 : OAI222_X1 port map( A1 => n2390, A2 => n769, B1 => n2422, B2 => n766
                           , C1 => n2358, C2 => n763, ZN => n3802);
   U3271 : NOR4_X1 port map( A1 => n5194, A2 => n5195, A3 => n5196, A4 => n5197
                           , ZN => n5193);
   U3272 : OAI22_X1 port map( A1 => n1845, A2 => n490, B1 => n1877, B2 => n487,
                           ZN => n5197);
   U3273 : OAI222_X1 port map( A1 => n2133, A2 => n466, B1 => n2165_port, B2 =>
                           n463, C1 => n2101, C2 => n460, ZN => n5194);
   U3274 : OAI222_X1 port map( A1 => n2037, A2 => n475, B1 => n2069, B2 => n472
                           , C1 => n2005, C2 => n469, ZN => n5195);
   U3275 : NOR4_X1 port map( A1 => n5203, A2 => n5204, A3 => n5205, A4 => n5206
                           , ZN => n5202);
   U3276 : OAI22_X1 port map( A1 => n2197, A2 => n72, B1 => n2229, B2 => n69, 
                           ZN => n5206);
   U3277 : OAI222_X1 port map( A1 => n2485, A2 => n48, B1 => n2517, B2 => n45, 
                           C1 => n2453, C2 => n42, ZN => n5203);
   U3278 : OAI222_X1 port map( A1 => n2389, A2 => n57, B1 => n2421, B2 => n54, 
                           C1 => n2357, C2 => n51, ZN => n5204);
   U3279 : NOR4_X1 port map( A1 => n3751, A2 => n3752, A3 => n3753, A4 => n3754
                           , ZN => n3750);
   U3280 : OAI22_X1 port map( A1 => n1845, A2 => n1298, B1 => n1877, B2 => 
                           n1199, ZN => n3754);
   U3281 : OAI222_X1 port map( A1 => n2133, A2 => n1178, B1 => n2165_port, B2 
                           => n1175, C1 => n2101, C2 => n1172, ZN => n3751);
   U3282 : OAI222_X1 port map( A1 => n2037, A2 => n1187, B1 => n2069, B2 => 
                           n1184, C1 => n2005, C2 => n1181, ZN => n3752);
   U3283 : NOR4_X1 port map( A1 => n3760, A2 => n3761, A3 => n3762, A4 => n3763
                           , ZN => n3759);
   U3284 : OAI22_X1 port map( A1 => n2197, A2 => n1136, B1 => n2229, B2 => n781
                           , ZN => n3763);
   U3285 : OAI222_X1 port map( A1 => n2485, A2 => n760, B1 => n2517, B2 => n757
                           , C1 => n2453, C2 => n754, ZN => n3760);
   U3286 : OAI222_X1 port map( A1 => n2389, A2 => n769, B1 => n2421, B2 => n766
                           , C1 => n2357, C2 => n763, ZN => n3761);
   U3287 : NOR4_X1 port map( A1 => n5153, A2 => n5154, A3 => n5155, A4 => n5156
                           , ZN => n5152);
   U3288 : OAI22_X1 port map( A1 => n1844, A2 => n490, B1 => n1876, B2 => n487,
                           ZN => n5156);
   U3289 : OAI222_X1 port map( A1 => n2132, A2 => n466, B1 => n2164_port, B2 =>
                           n463, C1 => n2100, C2 => n460, ZN => n5153);
   U3290 : OAI222_X1 port map( A1 => n2036, A2 => n475, B1 => n2068, B2 => n472
                           , C1 => n2004, C2 => n469, ZN => n5154);
   U3291 : NOR4_X1 port map( A1 => n5162, A2 => n5163, A3 => n5164, A4 => n5165
                           , ZN => n5161);
   U3292 : OAI22_X1 port map( A1 => n2196, A2 => n72, B1 => n2228, B2 => n69, 
                           ZN => n5165);
   U3293 : OAI222_X1 port map( A1 => n2484, A2 => n48, B1 => n2516, B2 => n45, 
                           C1 => n2452, C2 => n42, ZN => n5162);
   U3294 : OAI222_X1 port map( A1 => n2388, A2 => n57, B1 => n2420, B2 => n54, 
                           C1 => n2356, C2 => n51, ZN => n5163);
   U3295 : NOR4_X1 port map( A1 => n3710, A2 => n3711, A3 => n3712, A4 => n3713
                           , ZN => n3709);
   U3296 : OAI22_X1 port map( A1 => n1844, A2 => n1298, B1 => n1876, B2 => 
                           n1199, ZN => n3713);
   U3297 : OAI222_X1 port map( A1 => n2132, A2 => n1178, B1 => n2164_port, B2 
                           => n1175, C1 => n2100, C2 => n1172, ZN => n3710);
   U3298 : OAI222_X1 port map( A1 => n2036, A2 => n1187, B1 => n2068, B2 => 
                           n1184, C1 => n2004, C2 => n1181, ZN => n3711);
   U3299 : NOR4_X1 port map( A1 => n3719, A2 => n3720, A3 => n3721, A4 => n3722
                           , ZN => n3718);
   U3300 : OAI22_X1 port map( A1 => n2196, A2 => n1136, B1 => n2228, B2 => n781
                           , ZN => n3722);
   U3301 : OAI222_X1 port map( A1 => n2484, A2 => n760, B1 => n2516, B2 => n757
                           , C1 => n2452, C2 => n754, ZN => n3719);
   U3302 : OAI222_X1 port map( A1 => n2388, A2 => n769, B1 => n2420, B2 => n766
                           , C1 => n2356, C2 => n763, ZN => n3720);
   U3303 : NOR4_X1 port map( A1 => n5112, A2 => n5113, A3 => n5114, A4 => n5115
                           , ZN => n5111);
   U3304 : OAI22_X1 port map( A1 => n1843, A2 => n490, B1 => n1875, B2 => n487,
                           ZN => n5115);
   U3305 : OAI222_X1 port map( A1 => n2131, A2 => n466, B1 => n2163_port, B2 =>
                           n463, C1 => n2099, C2 => n460, ZN => n5112);
   U3306 : OAI222_X1 port map( A1 => n2035, A2 => n475, B1 => n2067, B2 => n472
                           , C1 => n2003, C2 => n469, ZN => n5113);
   U3307 : NOR4_X1 port map( A1 => n5121, A2 => n5122, A3 => n5123, A4 => n5124
                           , ZN => n5120);
   U3308 : OAI22_X1 port map( A1 => n2195, A2 => n72, B1 => n2227, B2 => n69, 
                           ZN => n5124);
   U3309 : OAI222_X1 port map( A1 => n2483, A2 => n48, B1 => n2515, B2 => n45, 
                           C1 => n2451, C2 => n42, ZN => n5121);
   U3310 : OAI222_X1 port map( A1 => n2387, A2 => n57, B1 => n2419, B2 => n54, 
                           C1 => n2355, C2 => n51, ZN => n5122);
   U3311 : NOR4_X1 port map( A1 => n3669, A2 => n3670, A3 => n3671, A4 => n3672
                           , ZN => n3668);
   U3312 : OAI22_X1 port map( A1 => n1843, A2 => n1298, B1 => n1875, B2 => 
                           n1199, ZN => n3672);
   U3313 : OAI222_X1 port map( A1 => n2131, A2 => n1178, B1 => n2163_port, B2 
                           => n1175, C1 => n2099, C2 => n1172, ZN => n3669);
   U3314 : OAI222_X1 port map( A1 => n2035, A2 => n1187, B1 => n2067, B2 => 
                           n1184, C1 => n2003, C2 => n1181, ZN => n3670);
   U3315 : NOR4_X1 port map( A1 => n3678, A2 => n3679, A3 => n3680, A4 => n3681
                           , ZN => n3677);
   U3316 : OAI22_X1 port map( A1 => n2195, A2 => n1136, B1 => n2227, B2 => n781
                           , ZN => n3681);
   U3317 : OAI222_X1 port map( A1 => n2483, A2 => n760, B1 => n2515, B2 => n757
                           , C1 => n2451, C2 => n754, ZN => n3678);
   U3318 : OAI222_X1 port map( A1 => n2387, A2 => n769, B1 => n2419, B2 => n766
                           , C1 => n2355, C2 => n763, ZN => n3679);
   U3319 : NOR4_X1 port map( A1 => n5071, A2 => n5072, A3 => n5073, A4 => n5074
                           , ZN => n5070);
   U3320 : OAI22_X1 port map( A1 => n1842, A2 => n490, B1 => n1874, B2 => n487,
                           ZN => n5074);
   U3321 : OAI222_X1 port map( A1 => n2130, A2 => n466, B1 => n2162, B2 => n463
                           , C1 => n2098, C2 => n460, ZN => n5071);
   U3322 : OAI222_X1 port map( A1 => n2034, A2 => n475, B1 => n2066, B2 => n472
                           , C1 => n2002, C2 => n469, ZN => n5072);
   U3323 : NOR4_X1 port map( A1 => n5080, A2 => n5081, A3 => n5082, A4 => n5083
                           , ZN => n5079);
   U3324 : OAI22_X1 port map( A1 => n2194, A2 => n72, B1 => n2226, B2 => n69, 
                           ZN => n5083);
   U3325 : OAI222_X1 port map( A1 => n2482, A2 => n48, B1 => n2514, B2 => n45, 
                           C1 => n2450, C2 => n42, ZN => n5080);
   U3326 : OAI222_X1 port map( A1 => n2386, A2 => n57, B1 => n2418, B2 => n54, 
                           C1 => n2354, C2 => n51, ZN => n5081);
   U3327 : NOR4_X1 port map( A1 => n3628, A2 => n3629, A3 => n3630, A4 => n3631
                           , ZN => n3627);
   U3328 : OAI22_X1 port map( A1 => n1842, A2 => n1298, B1 => n1874, B2 => 
                           n1199, ZN => n3631);
   U3329 : OAI222_X1 port map( A1 => n2130, A2 => n1178, B1 => n2162, B2 => 
                           n1175, C1 => n2098, C2 => n1172, ZN => n3628);
   U3330 : OAI222_X1 port map( A1 => n2034, A2 => n1187, B1 => n2066, B2 => 
                           n1184, C1 => n2002, C2 => n1181, ZN => n3629);
   U3331 : NOR4_X1 port map( A1 => n3637, A2 => n3638, A3 => n3639, A4 => n3640
                           , ZN => n3636);
   U3332 : OAI22_X1 port map( A1 => n2194, A2 => n1136, B1 => n2226, B2 => n781
                           , ZN => n3640);
   U3333 : OAI222_X1 port map( A1 => n2482, A2 => n760, B1 => n2514, B2 => n757
                           , C1 => n2450, C2 => n754, ZN => n3637);
   U3334 : OAI222_X1 port map( A1 => n2386, A2 => n769, B1 => n2418, B2 => n766
                           , C1 => n2354, C2 => n763, ZN => n3638);
   U3335 : NOR4_X1 port map( A1 => n5030, A2 => n5031, A3 => n5032, A4 => n5033
                           , ZN => n5029);
   U3336 : OAI22_X1 port map( A1 => n1841, A2 => n490, B1 => n1873, B2 => n487,
                           ZN => n5033);
   U3337 : OAI222_X1 port map( A1 => n2129, A2 => n466, B1 => n2161, B2 => n463
                           , C1 => n2097, C2 => n460, ZN => n5030);
   U3338 : OAI222_X1 port map( A1 => n2033, A2 => n475, B1 => n2065, B2 => n472
                           , C1 => n2001, C2 => n469, ZN => n5031);
   U3339 : NOR4_X1 port map( A1 => n5039, A2 => n5040, A3 => n5041, A4 => n5042
                           , ZN => n5038);
   U3340 : OAI22_X1 port map( A1 => n2193, A2 => n72, B1 => n2225, B2 => n69, 
                           ZN => n5042);
   U3341 : OAI222_X1 port map( A1 => n2481, A2 => n48, B1 => n2513, B2 => n45, 
                           C1 => n2449, C2 => n42, ZN => n5039);
   U3342 : OAI222_X1 port map( A1 => n2385, A2 => n57, B1 => n2417, B2 => n54, 
                           C1 => n2353, C2 => n51, ZN => n5040);
   U3343 : NOR4_X1 port map( A1 => n3587, A2 => n3588, A3 => n3589, A4 => n3590
                           , ZN => n3586);
   U3344 : OAI22_X1 port map( A1 => n1841, A2 => n1298, B1 => n1873, B2 => 
                           n1199, ZN => n3590);
   U3345 : OAI222_X1 port map( A1 => n2129, A2 => n1178, B1 => n2161, B2 => 
                           n1175, C1 => n2097, C2 => n1172, ZN => n3587);
   U3346 : OAI222_X1 port map( A1 => n2033, A2 => n1187, B1 => n2065, B2 => 
                           n1184, C1 => n2001, C2 => n1181, ZN => n3588);
   U3347 : NOR4_X1 port map( A1 => n3596, A2 => n3597, A3 => n3598, A4 => n3599
                           , ZN => n3595);
   U3348 : OAI22_X1 port map( A1 => n2193, A2 => n1136, B1 => n2225, B2 => n781
                           , ZN => n3599);
   U3349 : OAI222_X1 port map( A1 => n2481, A2 => n760, B1 => n2513, B2 => n757
                           , C1 => n2449, C2 => n754, ZN => n3596);
   U3350 : OAI222_X1 port map( A1 => n2385, A2 => n769, B1 => n2417, B2 => n766
                           , C1 => n2353, C2 => n763, ZN => n3597);
   U3351 : NOR4_X1 port map( A1 => n4945, A2 => n4946, A3 => n4947, A4 => n4948
                           , ZN => n4944);
   U3352 : OAI22_X1 port map( A1 => n1840, A2 => n490, B1 => n1872, B2 => n487,
                           ZN => n4948);
   U3353 : OAI222_X1 port map( A1 => n2128, A2 => n466, B1 => n2160, B2 => n463
                           , C1 => n2096, C2 => n460, ZN => n4945);
   U3354 : OAI222_X1 port map( A1 => n2032, A2 => n475, B1 => n2064, B2 => n472
                           , C1 => n2000, C2 => n469, ZN => n4946);
   U3355 : NOR4_X1 port map( A1 => n4976, A2 => n4977, A3 => n4978, A4 => n4979
                           , ZN => n4975);
   U3356 : OAI22_X1 port map( A1 => n2192, A2 => n72, B1 => n2224, B2 => n69, 
                           ZN => n4979);
   U3357 : OAI222_X1 port map( A1 => n2480, A2 => n48, B1 => n2512, B2 => n45, 
                           C1 => n2448, C2 => n42, ZN => n4976);
   U3358 : OAI222_X1 port map( A1 => n2384, A2 => n57, B1 => n2416, B2 => n54, 
                           C1 => n2352, C2 => n51, ZN => n4977);
   U3359 : NOR4_X1 port map( A1 => n3502, A2 => n3503, A3 => n3504, A4 => n3505
                           , ZN => n3501);
   U3360 : OAI22_X1 port map( A1 => n1840, A2 => n1298, B1 => n1872, B2 => 
                           n1199, ZN => n3505);
   U3361 : OAI222_X1 port map( A1 => n2128, A2 => n1178, B1 => n2160, B2 => 
                           n1175, C1 => n2096, C2 => n1172, ZN => n3502);
   U3362 : OAI222_X1 port map( A1 => n2032, A2 => n1187, B1 => n2064, B2 => 
                           n1184, C1 => n2000, C2 => n1181, ZN => n3503);
   U3363 : NOR4_X1 port map( A1 => n3533, A2 => n3534, A3 => n3535, A4 => n3536
                           , ZN => n3532);
   U3364 : OAI22_X1 port map( A1 => n2192, A2 => n1136, B1 => n2224, B2 => n781
                           , ZN => n3536);
   U3365 : OAI222_X1 port map( A1 => n2480, A2 => n760, B1 => n2512, B2 => n757
                           , C1 => n2448, C2 => n754, ZN => n3533);
   U3366 : OAI222_X1 port map( A1 => n2384, A2 => n769, B1 => n2416, B2 => n766
                           , C1 => n2352, C2 => n763, ZN => n3534);
   U3367 : AOI22_X1 port map( A1 => ADD_WR(1), A2 => n3391, B1 => N2154, B2 => 
                           N2151, ZN => n3406);
   U3368 : AOI22_X1 port map( A1 => N2163, A2 => n3391, B1 => N2156, B2 => 
                           N2151, ZN => n3359);
   U3369 : INV_X1 port map( A => ADD_WR(3), ZN => N2163);
   U3370 : AOI22_X1 port map( A1 => ADD_WR(0), A2 => n3391, B1 => N2153, B2 => 
                           N2151, ZN => n3405);
   U3371 : AOI22_X1 port map( A1 => ADD_WR(2), A2 => n3391, B1 => N2155, B2 => 
                           N2151, ZN => n3377);
   U3372 : AOI221_X1 port map( B1 => n455, B2 => REGISTERS_45_0_port, C1 => 
                           n452, C2 => REGISTERS_44_0_port, A => n6299, ZN => 
                           n6290);
   U3373 : OAI222_X1 port map( A1 => n1615, A2 => n449, B1 => n1647, B2 => n446
                           , C1 => n1583, C2 => n443, ZN => n6299);
   U3374 : AOI221_X1 port map( B1 => n37, B2 => REGISTERS_78_0_port, C1 => n34,
                           C2 => REGISTERS_77_0_port, A => n6311, ZN => n6303);
   U3375 : OAI222_X1 port map( A1 => n2671, A2 => n31, B1 => n2703, B2 => n28, 
                           C1 => n2639, C2 => n25, ZN => n6311);
   U3376 : AOI221_X1 port map( B1 => n1167, B2 => REGISTERS_45_0_port, C1 => 
                           n1164, C2 => REGISTERS_44_0_port, A => n4856, ZN => 
                           n4847);
   U3377 : OAI222_X1 port map( A1 => n1615, A2 => n1161, B1 => n1647, B2 => 
                           n1158, C1 => n1583, C2 => n1155, ZN => n4856);
   U3378 : AOI221_X1 port map( B1 => n749, B2 => REGISTERS_78_0_port, C1 => 
                           n746, C2 => REGISTERS_77_0_port, A => n4868, ZN => 
                           n4860);
   U3379 : OAI222_X1 port map( A1 => n2671, A2 => n743, B1 => n2703, B2 => n740
                           , C1 => n2639, C2 => n737, ZN => n4868);
   U3380 : AOI221_X1 port map( B1 => n455, B2 => REGISTERS_45_1_port, C1 => 
                           n452, C2 => REGISTERS_44_1_port, A => n6223, ZN => 
                           n6217);
   U3381 : OAI222_X1 port map( A1 => n1614, A2 => n449, B1 => n1646, B2 => n446
                           , C1 => n1582, C2 => n443, ZN => n6223);
   U3382 : AOI221_X1 port map( B1 => n37, B2 => REGISTERS_78_1_port, C1 => n34,
                           C2 => REGISTERS_77_1_port, A => n6232, ZN => n6226);
   U3383 : OAI222_X1 port map( A1 => n2670, A2 => n31, B1 => n2702, B2 => n28, 
                           C1 => n2638, C2 => n25, ZN => n6232);
   U3384 : AOI221_X1 port map( B1 => n1167, B2 => REGISTERS_45_1_port, C1 => 
                           n1164, C2 => REGISTERS_44_1_port, A => n4780, ZN => 
                           n4774);
   U3385 : OAI222_X1 port map( A1 => n1614, A2 => n1161, B1 => n1646, B2 => 
                           n1158, C1 => n1582, C2 => n1155, ZN => n4780);
   U3386 : AOI221_X1 port map( B1 => n749, B2 => REGISTERS_78_1_port, C1 => 
                           n746, C2 => REGISTERS_77_1_port, A => n4789, ZN => 
                           n4783);
   U3387 : OAI222_X1 port map( A1 => n2670, A2 => n743, B1 => n2702, B2 => n740
                           , C1 => n2638, C2 => n737, ZN => n4789);
   U3388 : AOI221_X1 port map( B1 => n455, B2 => REGISTERS_45_2_port, C1 => 
                           n452, C2 => REGISTERS_44_2_port, A => n6182, ZN => 
                           n6176);
   U3389 : OAI222_X1 port map( A1 => n1613, A2 => n449, B1 => n1645, B2 => n446
                           , C1 => n1581, C2 => n443, ZN => n6182);
   U3390 : AOI221_X1 port map( B1 => n37, B2 => REGISTERS_78_2_port, C1 => n34,
                           C2 => REGISTERS_77_2_port, A => n6191, ZN => n6185);
   U3391 : OAI222_X1 port map( A1 => n2669, A2 => n31, B1 => n2701, B2 => n28, 
                           C1 => n2637, C2 => n25, ZN => n6191);
   U3392 : AOI221_X1 port map( B1 => n1167, B2 => REGISTERS_45_2_port, C1 => 
                           n1164, C2 => REGISTERS_44_2_port, A => n4739, ZN => 
                           n4733);
   U3393 : OAI222_X1 port map( A1 => n1613, A2 => n1161, B1 => n1645, B2 => 
                           n1158, C1 => n1581, C2 => n1155, ZN => n4739);
   U3394 : AOI221_X1 port map( B1 => n749, B2 => REGISTERS_78_2_port, C1 => 
                           n746, C2 => REGISTERS_77_2_port, A => n4748, ZN => 
                           n4742);
   U3395 : OAI222_X1 port map( A1 => n2669, A2 => n743, B1 => n2701, B2 => n740
                           , C1 => n2637, C2 => n737, ZN => n4748);
   U3396 : AOI221_X1 port map( B1 => n455, B2 => REGISTERS_45_3_port, C1 => 
                           n452, C2 => REGISTERS_44_3_port, A => n6141, ZN => 
                           n6135);
   U3397 : OAI222_X1 port map( A1 => n1612, A2 => n449, B1 => n1644, B2 => n446
                           , C1 => n1580, C2 => n443, ZN => n6141);
   U3398 : AOI221_X1 port map( B1 => n37, B2 => REGISTERS_78_3_port, C1 => n34,
                           C2 => REGISTERS_77_3_port, A => n6150, ZN => n6144);
   U3399 : OAI222_X1 port map( A1 => n2668, A2 => n31, B1 => n2700, B2 => n28, 
                           C1 => n2636, C2 => n25, ZN => n6150);
   U3400 : AOI221_X1 port map( B1 => n1167, B2 => REGISTERS_45_3_port, C1 => 
                           n1164, C2 => REGISTERS_44_3_port, A => n4698, ZN => 
                           n4692);
   U3401 : OAI222_X1 port map( A1 => n1612, A2 => n1161, B1 => n1644, B2 => 
                           n1158, C1 => n1580, C2 => n1155, ZN => n4698);
   U3402 : AOI221_X1 port map( B1 => n749, B2 => REGISTERS_78_3_port, C1 => 
                           n746, C2 => REGISTERS_77_3_port, A => n4707, ZN => 
                           n4701);
   U3403 : OAI222_X1 port map( A1 => n2668, A2 => n743, B1 => n2700, B2 => n740
                           , C1 => n2636, C2 => n737, ZN => n4707);
   U3404 : AOI221_X1 port map( B1 => n455, B2 => REGISTERS_45_4_port, C1 => 
                           n452, C2 => REGISTERS_44_4_port, A => n6100, ZN => 
                           n6094);
   U3405 : OAI222_X1 port map( A1 => n1611, A2 => n449, B1 => n1643, B2 => n446
                           , C1 => n1579, C2 => n443, ZN => n6100);
   U3406 : AOI221_X1 port map( B1 => n37, B2 => REGISTERS_78_4_port, C1 => n34,
                           C2 => REGISTERS_77_4_port, A => n6109, ZN => n6103);
   U3407 : OAI222_X1 port map( A1 => n2667, A2 => n31, B1 => n2699, B2 => n28, 
                           C1 => n2635, C2 => n25, ZN => n6109);
   U3408 : AOI221_X1 port map( B1 => n1167, B2 => REGISTERS_45_4_port, C1 => 
                           n1164, C2 => REGISTERS_44_4_port, A => n4657, ZN => 
                           n4651);
   U3409 : OAI222_X1 port map( A1 => n1611, A2 => n1161, B1 => n1643, B2 => 
                           n1158, C1 => n1579, C2 => n1155, ZN => n4657);
   U3410 : AOI221_X1 port map( B1 => n749, B2 => REGISTERS_78_4_port, C1 => 
                           n746, C2 => REGISTERS_77_4_port, A => n4666, ZN => 
                           n4660);
   U3411 : OAI222_X1 port map( A1 => n2667, A2 => n743, B1 => n2699, B2 => n740
                           , C1 => n2635, C2 => n737, ZN => n4666);
   U3412 : AOI221_X1 port map( B1 => n455, B2 => REGISTERS_45_5_port, C1 => 
                           n452, C2 => REGISTERS_44_5_port, A => n6059, ZN => 
                           n6053);
   U3413 : OAI222_X1 port map( A1 => n1610, A2 => n449, B1 => n1642, B2 => n446
                           , C1 => n1578, C2 => n443, ZN => n6059);
   U3414 : AOI221_X1 port map( B1 => n37, B2 => REGISTERS_78_5_port, C1 => n34,
                           C2 => REGISTERS_77_5_port, A => n6068, ZN => n6062);
   U3415 : OAI222_X1 port map( A1 => n2666, A2 => n31, B1 => n2698, B2 => n28, 
                           C1 => n2634, C2 => n25, ZN => n6068);
   U3416 : AOI221_X1 port map( B1 => n1167, B2 => REGISTERS_45_5_port, C1 => 
                           n1164, C2 => REGISTERS_44_5_port, A => n4616, ZN => 
                           n4610);
   U3417 : OAI222_X1 port map( A1 => n1610, A2 => n1161, B1 => n1642, B2 => 
                           n1158, C1 => n1578, C2 => n1155, ZN => n4616);
   U3418 : AOI221_X1 port map( B1 => n749, B2 => REGISTERS_78_5_port, C1 => 
                           n746, C2 => REGISTERS_77_5_port, A => n4625, ZN => 
                           n4619);
   U3419 : OAI222_X1 port map( A1 => n2666, A2 => n743, B1 => n2698, B2 => n740
                           , C1 => n2634, C2 => n737, ZN => n4625);
   U3420 : AOI221_X1 port map( B1 => n455, B2 => REGISTERS_45_6_port, C1 => 
                           n452, C2 => REGISTERS_44_6_port, A => n6018, ZN => 
                           n6012);
   U3421 : OAI222_X1 port map( A1 => n1609, A2 => n449, B1 => n1641, B2 => n446
                           , C1 => n1577, C2 => n443, ZN => n6018);
   U3422 : AOI221_X1 port map( B1 => n37, B2 => REGISTERS_78_6_port, C1 => n34,
                           C2 => REGISTERS_77_6_port, A => n6027, ZN => n6021);
   U3423 : OAI222_X1 port map( A1 => n2665, A2 => n31, B1 => n2697, B2 => n28, 
                           C1 => n2633, C2 => n25, ZN => n6027);
   U3424 : AOI221_X1 port map( B1 => n1167, B2 => REGISTERS_45_6_port, C1 => 
                           n1164, C2 => REGISTERS_44_6_port, A => n4575, ZN => 
                           n4569);
   U3425 : OAI222_X1 port map( A1 => n1609, A2 => n1161, B1 => n1641, B2 => 
                           n1158, C1 => n1577, C2 => n1155, ZN => n4575);
   U3426 : AOI221_X1 port map( B1 => n749, B2 => REGISTERS_78_6_port, C1 => 
                           n746, C2 => REGISTERS_77_6_port, A => n4584, ZN => 
                           n4578);
   U3427 : OAI222_X1 port map( A1 => n2665, A2 => n743, B1 => n2697, B2 => n740
                           , C1 => n2633, C2 => n737, ZN => n4584);
   U3428 : AOI221_X1 port map( B1 => n455, B2 => REGISTERS_45_7_port, C1 => 
                           n452, C2 => REGISTERS_44_7_port, A => n5977, ZN => 
                           n5971);
   U3429 : OAI222_X1 port map( A1 => n1608, A2 => n449, B1 => n1640, B2 => n446
                           , C1 => n1576, C2 => n443, ZN => n5977);
   U3430 : AOI221_X1 port map( B1 => n37, B2 => REGISTERS_78_7_port, C1 => n34,
                           C2 => REGISTERS_77_7_port, A => n5986, ZN => n5980);
   U3431 : OAI222_X1 port map( A1 => n2664, A2 => n31, B1 => n2696, B2 => n28, 
                           C1 => n2632, C2 => n25, ZN => n5986);
   U3432 : AOI221_X1 port map( B1 => n1167, B2 => REGISTERS_45_7_port, C1 => 
                           n1164, C2 => REGISTERS_44_7_port, A => n4534, ZN => 
                           n4528);
   U3433 : OAI222_X1 port map( A1 => n1608, A2 => n1161, B1 => n1640, B2 => 
                           n1158, C1 => n1576, C2 => n1155, ZN => n4534);
   U3434 : AOI221_X1 port map( B1 => n749, B2 => REGISTERS_78_7_port, C1 => 
                           n746, C2 => REGISTERS_77_7_port, A => n4543, ZN => 
                           n4537);
   U3435 : OAI222_X1 port map( A1 => n2664, A2 => n743, B1 => n2696, B2 => n740
                           , C1 => n2632, C2 => n737, ZN => n4543);
   U3436 : AOI221_X1 port map( B1 => n455, B2 => REGISTERS_45_8_port, C1 => 
                           n452, C2 => REGISTERS_44_8_port, A => n5936, ZN => 
                           n5930);
   U3437 : OAI222_X1 port map( A1 => n1607, A2 => n449, B1 => n1639, B2 => n446
                           , C1 => n1575, C2 => n443, ZN => n5936);
   U3438 : AOI221_X1 port map( B1 => n37, B2 => REGISTERS_78_8_port, C1 => n34,
                           C2 => REGISTERS_77_8_port, A => n5945, ZN => n5939);
   U3439 : OAI222_X1 port map( A1 => n2663, A2 => n31, B1 => n2695, B2 => n28, 
                           C1 => n2631, C2 => n25, ZN => n5945);
   U3440 : AOI221_X1 port map( B1 => n1167, B2 => REGISTERS_45_8_port, C1 => 
                           n1164, C2 => REGISTERS_44_8_port, A => n4493, ZN => 
                           n4487);
   U3441 : OAI222_X1 port map( A1 => n1607, A2 => n1161, B1 => n1639, B2 => 
                           n1158, C1 => n1575, C2 => n1155, ZN => n4493);
   U3442 : AOI221_X1 port map( B1 => n749, B2 => REGISTERS_78_8_port, C1 => 
                           n746, C2 => REGISTERS_77_8_port, A => n4502, ZN => 
                           n4496);
   U3443 : OAI222_X1 port map( A1 => n2663, A2 => n743, B1 => n2695, B2 => n740
                           , C1 => n2631, C2 => n737, ZN => n4502);
   U3444 : AOI221_X1 port map( B1 => n455, B2 => REGISTERS_45_9_port, C1 => 
                           n452, C2 => REGISTERS_44_9_port, A => n5895, ZN => 
                           n5889);
   U3445 : OAI222_X1 port map( A1 => n1606, A2 => n449, B1 => n1638, B2 => n446
                           , C1 => n1574, C2 => n443, ZN => n5895);
   U3446 : AOI221_X1 port map( B1 => n37, B2 => REGISTERS_78_9_port, C1 => n34,
                           C2 => REGISTERS_77_9_port, A => n5904, ZN => n5898);
   U3447 : OAI222_X1 port map( A1 => n2662, A2 => n31, B1 => n2694, B2 => n28, 
                           C1 => n2630, C2 => n25, ZN => n5904);
   U3448 : AOI221_X1 port map( B1 => n1167, B2 => REGISTERS_45_9_port, C1 => 
                           n1164, C2 => REGISTERS_44_9_port, A => n4452, ZN => 
                           n4446);
   U3449 : OAI222_X1 port map( A1 => n1606, A2 => n1161, B1 => n1638, B2 => 
                           n1158, C1 => n1574, C2 => n1155, ZN => n4452);
   U3450 : AOI221_X1 port map( B1 => n749, B2 => REGISTERS_78_9_port, C1 => 
                           n746, C2 => REGISTERS_77_9_port, A => n4461, ZN => 
                           n4455);
   U3451 : OAI222_X1 port map( A1 => n2662, A2 => n743, B1 => n2694, B2 => n740
                           , C1 => n2630, C2 => n737, ZN => n4461);
   U3452 : AOI221_X1 port map( B1 => n455, B2 => REGISTERS_45_10_port, C1 => 
                           n452, C2 => REGISTERS_44_10_port, A => n5854, ZN => 
                           n5848);
   U3453 : OAI222_X1 port map( A1 => n1605, A2 => n449, B1 => n1637, B2 => n446
                           , C1 => n1573, C2 => n443, ZN => n5854);
   U3454 : AOI221_X1 port map( B1 => n37, B2 => REGISTERS_78_10_port, C1 => n34
                           , C2 => REGISTERS_77_10_port, A => n5863, ZN => 
                           n5857);
   U3455 : OAI222_X1 port map( A1 => n2661, A2 => n31, B1 => n2693, B2 => n28, 
                           C1 => n2629, C2 => n25, ZN => n5863);
   U3456 : AOI221_X1 port map( B1 => n1167, B2 => REGISTERS_45_10_port, C1 => 
                           n1164, C2 => REGISTERS_44_10_port, A => n4411, ZN =>
                           n4405);
   U3457 : OAI222_X1 port map( A1 => n1605, A2 => n1161, B1 => n1637, B2 => 
                           n1158, C1 => n1573, C2 => n1155, ZN => n4411);
   U3458 : AOI221_X1 port map( B1 => n749, B2 => REGISTERS_78_10_port, C1 => 
                           n746, C2 => REGISTERS_77_10_port, A => n4420, ZN => 
                           n4414);
   U3459 : OAI222_X1 port map( A1 => n2661, A2 => n743, B1 => n2693, B2 => n740
                           , C1 => n2629, C2 => n737, ZN => n4420);
   U3460 : AOI221_X1 port map( B1 => n455, B2 => REGISTERS_45_11_port, C1 => 
                           n452, C2 => REGISTERS_44_11_port, A => n5813, ZN => 
                           n5807);
   U3461 : OAI222_X1 port map( A1 => n1604, A2 => n449, B1 => n1636, B2 => n446
                           , C1 => n1572, C2 => n443, ZN => n5813);
   U3462 : AOI221_X1 port map( B1 => n37, B2 => REGISTERS_78_11_port, C1 => n34
                           , C2 => REGISTERS_77_11_port, A => n5822, ZN => 
                           n5816);
   U3463 : OAI222_X1 port map( A1 => n2660, A2 => n31, B1 => n2692, B2 => n28, 
                           C1 => n2628, C2 => n25, ZN => n5822);
   U3464 : AOI221_X1 port map( B1 => n1167, B2 => REGISTERS_45_11_port, C1 => 
                           n1164, C2 => REGISTERS_44_11_port, A => n4370, ZN =>
                           n4364);
   U3465 : OAI222_X1 port map( A1 => n1604, A2 => n1161, B1 => n1636, B2 => 
                           n1158, C1 => n1572, C2 => n1155, ZN => n4370);
   U3466 : AOI221_X1 port map( B1 => n749, B2 => REGISTERS_78_11_port, C1 => 
                           n746, C2 => REGISTERS_77_11_port, A => n4379, ZN => 
                           n4373);
   U3467 : OAI222_X1 port map( A1 => n2660, A2 => n743, B1 => n2692, B2 => n740
                           , C1 => n2628, C2 => n737, ZN => n4379);
   U3468 : AOI221_X1 port map( B1 => n456, B2 => REGISTERS_45_12_port, C1 => 
                           n453, C2 => REGISTERS_44_12_port, A => n5772, ZN => 
                           n5766);
   U3469 : OAI222_X1 port map( A1 => n1603, A2 => n450, B1 => n1635, B2 => n447
                           , C1 => n1571, C2 => n444, ZN => n5772);
   U3470 : AOI221_X1 port map( B1 => n38, B2 => REGISTERS_78_12_port, C1 => n35
                           , C2 => REGISTERS_77_12_port, A => n5781, ZN => 
                           n5775);
   U3471 : OAI222_X1 port map( A1 => n2659, A2 => n32, B1 => n2691, B2 => n29, 
                           C1 => n2627, C2 => n26, ZN => n5781);
   U3472 : AOI221_X1 port map( B1 => n1168, B2 => REGISTERS_45_12_port, C1 => 
                           n1165, C2 => REGISTERS_44_12_port, A => n4329, ZN =>
                           n4323);
   U3473 : OAI222_X1 port map( A1 => n1603, A2 => n1162, B1 => n1635, B2 => 
                           n1159, C1 => n1571, C2 => n1156, ZN => n4329);
   U3474 : AOI221_X1 port map( B1 => n750, B2 => REGISTERS_78_12_port, C1 => 
                           n747, C2 => REGISTERS_77_12_port, A => n4338, ZN => 
                           n4332);
   U3475 : OAI222_X1 port map( A1 => n2659, A2 => n744, B1 => n2691, B2 => n741
                           , C1 => n2627, C2 => n738, ZN => n4338);
   U3476 : AOI221_X1 port map( B1 => n456, B2 => REGISTERS_45_13_port, C1 => 
                           n453, C2 => REGISTERS_44_13_port, A => n5731, ZN => 
                           n5725);
   U3477 : OAI222_X1 port map( A1 => n1602, A2 => n450, B1 => n1634, B2 => n447
                           , C1 => n1570, C2 => n444, ZN => n5731);
   U3478 : AOI221_X1 port map( B1 => n38, B2 => REGISTERS_78_13_port, C1 => n35
                           , C2 => REGISTERS_77_13_port, A => n5740, ZN => 
                           n5734);
   U3479 : OAI222_X1 port map( A1 => n2658, A2 => n32, B1 => n2690, B2 => n29, 
                           C1 => n2626, C2 => n26, ZN => n5740);
   U3480 : AOI221_X1 port map( B1 => n1168, B2 => REGISTERS_45_13_port, C1 => 
                           n1165, C2 => REGISTERS_44_13_port, A => n4288, ZN =>
                           n4282);
   U3481 : OAI222_X1 port map( A1 => n1602, A2 => n1162, B1 => n1634, B2 => 
                           n1159, C1 => n1570, C2 => n1156, ZN => n4288);
   U3482 : AOI221_X1 port map( B1 => n750, B2 => REGISTERS_78_13_port, C1 => 
                           n747, C2 => REGISTERS_77_13_port, A => n4297, ZN => 
                           n4291);
   U3483 : OAI222_X1 port map( A1 => n2658, A2 => n744, B1 => n2690, B2 => n741
                           , C1 => n2626, C2 => n738, ZN => n4297);
   U3484 : AOI221_X1 port map( B1 => n456, B2 => REGISTERS_45_14_port, C1 => 
                           n453, C2 => REGISTERS_44_14_port, A => n5690, ZN => 
                           n5684);
   U3485 : OAI222_X1 port map( A1 => n1601, A2 => n450, B1 => n1633, B2 => n447
                           , C1 => n1569, C2 => n444, ZN => n5690);
   U3486 : AOI221_X1 port map( B1 => n38, B2 => REGISTERS_78_14_port, C1 => n35
                           , C2 => REGISTERS_77_14_port, A => n5699, ZN => 
                           n5693);
   U3487 : OAI222_X1 port map( A1 => n2657, A2 => n32, B1 => n2689, B2 => n29, 
                           C1 => n2625, C2 => n26, ZN => n5699);
   U3488 : AOI221_X1 port map( B1 => n1168, B2 => REGISTERS_45_14_port, C1 => 
                           n1165, C2 => REGISTERS_44_14_port, A => n4247, ZN =>
                           n4241);
   U3489 : OAI222_X1 port map( A1 => n1601, A2 => n1162, B1 => n1633, B2 => 
                           n1159, C1 => n1569, C2 => n1156, ZN => n4247);
   U3490 : AOI221_X1 port map( B1 => n750, B2 => REGISTERS_78_14_port, C1 => 
                           n747, C2 => REGISTERS_77_14_port, A => n4256, ZN => 
                           n4250);
   U3491 : OAI222_X1 port map( A1 => n2657, A2 => n744, B1 => n2689, B2 => n741
                           , C1 => n2625, C2 => n738, ZN => n4256);
   U3492 : AOI221_X1 port map( B1 => n456, B2 => REGISTERS_45_15_port, C1 => 
                           n453, C2 => REGISTERS_44_15_port, A => n5649, ZN => 
                           n5643);
   U3493 : OAI222_X1 port map( A1 => n1600, A2 => n450, B1 => n1632, B2 => n447
                           , C1 => n1568, C2 => n444, ZN => n5649);
   U3494 : AOI221_X1 port map( B1 => n38, B2 => REGISTERS_78_15_port, C1 => n35
                           , C2 => REGISTERS_77_15_port, A => n5658, ZN => 
                           n5652);
   U3495 : OAI222_X1 port map( A1 => n2656, A2 => n32, B1 => n2688, B2 => n29, 
                           C1 => n2624, C2 => n26, ZN => n5658);
   U3496 : AOI221_X1 port map( B1 => n1168, B2 => REGISTERS_45_15_port, C1 => 
                           n1165, C2 => REGISTERS_44_15_port, A => n4206, ZN =>
                           n4200);
   U3497 : OAI222_X1 port map( A1 => n1600, A2 => n1162, B1 => n1632, B2 => 
                           n1159, C1 => n1568, C2 => n1156, ZN => n4206);
   U3498 : AOI221_X1 port map( B1 => n750, B2 => REGISTERS_78_15_port, C1 => 
                           n747, C2 => REGISTERS_77_15_port, A => n4215, ZN => 
                           n4209);
   U3499 : OAI222_X1 port map( A1 => n2656, A2 => n744, B1 => n2688, B2 => n741
                           , C1 => n2624, C2 => n738, ZN => n4215);
   U3500 : AOI221_X1 port map( B1 => n456, B2 => REGISTERS_45_16_port, C1 => 
                           n453, C2 => REGISTERS_44_16_port, A => n5608, ZN => 
                           n5602);
   U3501 : OAI222_X1 port map( A1 => n1599, A2 => n450, B1 => n1631, B2 => n447
                           , C1 => n1567, C2 => n444, ZN => n5608);
   U3502 : AOI221_X1 port map( B1 => n38, B2 => REGISTERS_78_16_port, C1 => n35
                           , C2 => REGISTERS_77_16_port, A => n5617, ZN => 
                           n5611);
   U3503 : OAI222_X1 port map( A1 => n2655, A2 => n32, B1 => n2687, B2 => n29, 
                           C1 => n2623, C2 => n26, ZN => n5617);
   U3504 : AOI221_X1 port map( B1 => n1168, B2 => REGISTERS_45_16_port, C1 => 
                           n1165, C2 => REGISTERS_44_16_port, A => n4165, ZN =>
                           n4159);
   U3505 : OAI222_X1 port map( A1 => n1599, A2 => n1162, B1 => n1631, B2 => 
                           n1159, C1 => n1567, C2 => n1156, ZN => n4165);
   U3506 : AOI221_X1 port map( B1 => n750, B2 => REGISTERS_78_16_port, C1 => 
                           n747, C2 => REGISTERS_77_16_port, A => n4174, ZN => 
                           n4168);
   U3507 : OAI222_X1 port map( A1 => n2655, A2 => n744, B1 => n2687, B2 => n741
                           , C1 => n2623, C2 => n738, ZN => n4174);
   U3508 : AOI221_X1 port map( B1 => n456, B2 => REGISTERS_45_17_port, C1 => 
                           n453, C2 => REGISTERS_44_17_port, A => n5567, ZN => 
                           n5561);
   U3509 : OAI222_X1 port map( A1 => n1598, A2 => n450, B1 => n1630, B2 => n447
                           , C1 => n1566, C2 => n444, ZN => n5567);
   U3510 : AOI221_X1 port map( B1 => n38, B2 => REGISTERS_78_17_port, C1 => n35
                           , C2 => REGISTERS_77_17_port, A => n5576, ZN => 
                           n5570);
   U3511 : OAI222_X1 port map( A1 => n2654, A2 => n32, B1 => n2686, B2 => n29, 
                           C1 => n2622, C2 => n26, ZN => n5576);
   U3512 : AOI221_X1 port map( B1 => n1168, B2 => REGISTERS_45_17_port, C1 => 
                           n1165, C2 => REGISTERS_44_17_port, A => n4124, ZN =>
                           n4118);
   U3513 : OAI222_X1 port map( A1 => n1598, A2 => n1162, B1 => n1630, B2 => 
                           n1159, C1 => n1566, C2 => n1156, ZN => n4124);
   U3514 : AOI221_X1 port map( B1 => n750, B2 => REGISTERS_78_17_port, C1 => 
                           n747, C2 => REGISTERS_77_17_port, A => n4133, ZN => 
                           n4127);
   U3515 : OAI222_X1 port map( A1 => n2654, A2 => n744, B1 => n2686, B2 => n741
                           , C1 => n2622, C2 => n738, ZN => n4133);
   U3516 : AOI221_X1 port map( B1 => n456, B2 => REGISTERS_45_18_port, C1 => 
                           n453, C2 => REGISTERS_44_18_port, A => n5526, ZN => 
                           n5520);
   U3517 : OAI222_X1 port map( A1 => n1597, A2 => n450, B1 => n1629, B2 => n447
                           , C1 => n1565, C2 => n444, ZN => n5526);
   U3518 : AOI221_X1 port map( B1 => n38, B2 => REGISTERS_78_18_port, C1 => n35
                           , C2 => REGISTERS_77_18_port, A => n5535, ZN => 
                           n5529);
   U3519 : OAI222_X1 port map( A1 => n2653, A2 => n32, B1 => n2685, B2 => n29, 
                           C1 => n2621, C2 => n26, ZN => n5535);
   U3520 : AOI221_X1 port map( B1 => n1168, B2 => REGISTERS_45_18_port, C1 => 
                           n1165, C2 => REGISTERS_44_18_port, A => n4083, ZN =>
                           n4077);
   U3521 : OAI222_X1 port map( A1 => n1597, A2 => n1162, B1 => n1629, B2 => 
                           n1159, C1 => n1565, C2 => n1156, ZN => n4083);
   U3522 : AOI221_X1 port map( B1 => n750, B2 => REGISTERS_78_18_port, C1 => 
                           n747, C2 => REGISTERS_77_18_port, A => n4092, ZN => 
                           n4086);
   U3523 : OAI222_X1 port map( A1 => n2653, A2 => n744, B1 => n2685, B2 => n741
                           , C1 => n2621, C2 => n738, ZN => n4092);
   U3524 : AOI221_X1 port map( B1 => n456, B2 => REGISTERS_45_19_port, C1 => 
                           n453, C2 => REGISTERS_44_19_port, A => n5485, ZN => 
                           n5479);
   U3525 : OAI222_X1 port map( A1 => n1596, A2 => n450, B1 => n1628, B2 => n447
                           , C1 => n1564, C2 => n444, ZN => n5485);
   U3526 : AOI221_X1 port map( B1 => n38, B2 => REGISTERS_78_19_port, C1 => n35
                           , C2 => REGISTERS_77_19_port, A => n5494, ZN => 
                           n5488);
   U3527 : OAI222_X1 port map( A1 => n2652, A2 => n32, B1 => n2684, B2 => n29, 
                           C1 => n2620, C2 => n26, ZN => n5494);
   U3528 : AOI221_X1 port map( B1 => n1168, B2 => REGISTERS_45_19_port, C1 => 
                           n1165, C2 => REGISTERS_44_19_port, A => n4042, ZN =>
                           n4036);
   U3529 : OAI222_X1 port map( A1 => n1596, A2 => n1162, B1 => n1628, B2 => 
                           n1159, C1 => n1564, C2 => n1156, ZN => n4042);
   U3530 : AOI221_X1 port map( B1 => n750, B2 => REGISTERS_78_19_port, C1 => 
                           n747, C2 => REGISTERS_77_19_port, A => n4051, ZN => 
                           n4045);
   U3531 : OAI222_X1 port map( A1 => n2652, A2 => n744, B1 => n2684, B2 => n741
                           , C1 => n2620, C2 => n738, ZN => n4051);
   U3532 : AOI221_X1 port map( B1 => n456, B2 => REGISTERS_45_20_port, C1 => 
                           n453, C2 => REGISTERS_44_20_port, A => n5444, ZN => 
                           n5438);
   U3533 : OAI222_X1 port map( A1 => n1595, A2 => n450, B1 => n1627, B2 => n447
                           , C1 => n1563, C2 => n444, ZN => n5444);
   U3534 : AOI221_X1 port map( B1 => n38, B2 => REGISTERS_78_20_port, C1 => n35
                           , C2 => REGISTERS_77_20_port, A => n5453, ZN => 
                           n5447);
   U3535 : OAI222_X1 port map( A1 => n2651, A2 => n32, B1 => n2683, B2 => n29, 
                           C1 => n2619, C2 => n26, ZN => n5453);
   U3536 : AOI221_X1 port map( B1 => n1168, B2 => REGISTERS_45_20_port, C1 => 
                           n1165, C2 => REGISTERS_44_20_port, A => n4001, ZN =>
                           n3995);
   U3537 : OAI222_X1 port map( A1 => n1595, A2 => n1162, B1 => n1627, B2 => 
                           n1159, C1 => n1563, C2 => n1156, ZN => n4001);
   U3538 : AOI221_X1 port map( B1 => n750, B2 => REGISTERS_78_20_port, C1 => 
                           n747, C2 => REGISTERS_77_20_port, A => n4010, ZN => 
                           n4004);
   U3539 : OAI222_X1 port map( A1 => n2651, A2 => n744, B1 => n2683, B2 => n741
                           , C1 => n2619, C2 => n738, ZN => n4010);
   U3540 : AOI221_X1 port map( B1 => n456, B2 => REGISTERS_45_21_port, C1 => 
                           n453, C2 => REGISTERS_44_21_port, A => n5403, ZN => 
                           n5397);
   U3541 : OAI222_X1 port map( A1 => n1594, A2 => n450, B1 => n1626, B2 => n447
                           , C1 => n1562, C2 => n444, ZN => n5403);
   U3542 : AOI221_X1 port map( B1 => n38, B2 => REGISTERS_78_21_port, C1 => n35
                           , C2 => REGISTERS_77_21_port, A => n5412, ZN => 
                           n5406);
   U3543 : OAI222_X1 port map( A1 => n2650, A2 => n32, B1 => n2682, B2 => n29, 
                           C1 => n2618, C2 => n26, ZN => n5412);
   U3544 : AOI221_X1 port map( B1 => n1168, B2 => REGISTERS_45_21_port, C1 => 
                           n1165, C2 => REGISTERS_44_21_port, A => n3960, ZN =>
                           n3954);
   U3545 : OAI222_X1 port map( A1 => n1594, A2 => n1162, B1 => n1626, B2 => 
                           n1159, C1 => n1562, C2 => n1156, ZN => n3960);
   U3546 : AOI221_X1 port map( B1 => n750, B2 => REGISTERS_78_21_port, C1 => 
                           n747, C2 => REGISTERS_77_21_port, A => n3969, ZN => 
                           n3963);
   U3547 : OAI222_X1 port map( A1 => n2650, A2 => n744, B1 => n2682, B2 => n741
                           , C1 => n2618, C2 => n738, ZN => n3969);
   U3548 : AOI221_X1 port map( B1 => n456, B2 => REGISTERS_45_22_port, C1 => 
                           n453, C2 => REGISTERS_44_22_port, A => n5362, ZN => 
                           n5356);
   U3549 : OAI222_X1 port map( A1 => n1593, A2 => n450, B1 => n1625, B2 => n447
                           , C1 => n1561, C2 => n444, ZN => n5362);
   U3550 : AOI221_X1 port map( B1 => n38, B2 => REGISTERS_78_22_port, C1 => n35
                           , C2 => REGISTERS_77_22_port, A => n5371, ZN => 
                           n5365);
   U3551 : OAI222_X1 port map( A1 => n2649, A2 => n32, B1 => n2681, B2 => n29, 
                           C1 => n2617, C2 => n26, ZN => n5371);
   U3552 : AOI221_X1 port map( B1 => n1168, B2 => REGISTERS_45_22_port, C1 => 
                           n1165, C2 => REGISTERS_44_22_port, A => n3919, ZN =>
                           n3913);
   U3553 : OAI222_X1 port map( A1 => n1593, A2 => n1162, B1 => n1625, B2 => 
                           n1159, C1 => n1561, C2 => n1156, ZN => n3919);
   U3554 : AOI221_X1 port map( B1 => n750, B2 => REGISTERS_78_22_port, C1 => 
                           n747, C2 => REGISTERS_77_22_port, A => n3928, ZN => 
                           n3922);
   U3555 : OAI222_X1 port map( A1 => n2649, A2 => n744, B1 => n2681, B2 => n741
                           , C1 => n2617, C2 => n738, ZN => n3928);
   U3556 : AOI221_X1 port map( B1 => n456, B2 => REGISTERS_45_23_port, C1 => 
                           n453, C2 => REGISTERS_44_23_port, A => n5321, ZN => 
                           n5315);
   U3557 : OAI222_X1 port map( A1 => n1592, A2 => n450, B1 => n1624, B2 => n447
                           , C1 => n1560, C2 => n444, ZN => n5321);
   U3558 : AOI221_X1 port map( B1 => n38, B2 => REGISTERS_78_23_port, C1 => n35
                           , C2 => REGISTERS_77_23_port, A => n5330, ZN => 
                           n5324);
   U3559 : OAI222_X1 port map( A1 => n2648, A2 => n32, B1 => n2680, B2 => n29, 
                           C1 => n2616, C2 => n26, ZN => n5330);
   U3560 : AOI221_X1 port map( B1 => n1168, B2 => REGISTERS_45_23_port, C1 => 
                           n1165, C2 => REGISTERS_44_23_port, A => n3878, ZN =>
                           n3872);
   U3561 : OAI222_X1 port map( A1 => n1592, A2 => n1162, B1 => n1624, B2 => 
                           n1159, C1 => n1560, C2 => n1156, ZN => n3878);
   U3562 : AOI221_X1 port map( B1 => n750, B2 => REGISTERS_78_23_port, C1 => 
                           n747, C2 => REGISTERS_77_23_port, A => n3887, ZN => 
                           n3881);
   U3563 : OAI222_X1 port map( A1 => n2648, A2 => n744, B1 => n2680, B2 => n741
                           , C1 => n2616, C2 => n738, ZN => n3887);
   U3564 : AOI221_X1 port map( B1 => n457, B2 => REGISTERS_45_24_port, C1 => 
                           n454, C2 => REGISTERS_44_24_port, A => n5280, ZN => 
                           n5274);
   U3565 : OAI222_X1 port map( A1 => n1591, A2 => n451, B1 => n1623, B2 => n448
                           , C1 => n1559, C2 => n445, ZN => n5280);
   U3566 : AOI221_X1 port map( B1 => n39, B2 => REGISTERS_78_24_port, C1 => n36
                           , C2 => REGISTERS_77_24_port, A => n5289, ZN => 
                           n5283);
   U3567 : OAI222_X1 port map( A1 => n2647, A2 => n33, B1 => n2679, B2 => n30, 
                           C1 => n2615, C2 => n27, ZN => n5289);
   U3568 : AOI221_X1 port map( B1 => n1169, B2 => REGISTERS_45_24_port, C1 => 
                           n1166, C2 => REGISTERS_44_24_port, A => n3837, ZN =>
                           n3831);
   U3569 : OAI222_X1 port map( A1 => n1591, A2 => n1163, B1 => n1623, B2 => 
                           n1160, C1 => n1559, C2 => n1157, ZN => n3837);
   U3570 : AOI221_X1 port map( B1 => n751, B2 => REGISTERS_78_24_port, C1 => 
                           n748, C2 => REGISTERS_77_24_port, A => n3846, ZN => 
                           n3840);
   U3571 : OAI222_X1 port map( A1 => n2647, A2 => n745, B1 => n2679, B2 => n742
                           , C1 => n2615, C2 => n739, ZN => n3846);
   U3572 : AOI221_X1 port map( B1 => n457, B2 => REGISTERS_45_25_port, C1 => 
                           n454, C2 => REGISTERS_44_25_port, A => n5239, ZN => 
                           n5233);
   U3573 : OAI222_X1 port map( A1 => n1590, A2 => n451, B1 => n1622, B2 => n448
                           , C1 => n1558, C2 => n445, ZN => n5239);
   U3574 : AOI221_X1 port map( B1 => n39, B2 => REGISTERS_78_25_port, C1 => n36
                           , C2 => REGISTERS_77_25_port, A => n5248, ZN => 
                           n5242);
   U3575 : OAI222_X1 port map( A1 => n2646, A2 => n33, B1 => n2678, B2 => n30, 
                           C1 => n2614, C2 => n27, ZN => n5248);
   U3576 : AOI221_X1 port map( B1 => n1169, B2 => REGISTERS_45_25_port, C1 => 
                           n1166, C2 => REGISTERS_44_25_port, A => n3796, ZN =>
                           n3790);
   U3577 : OAI222_X1 port map( A1 => n1590, A2 => n1163, B1 => n1622, B2 => 
                           n1160, C1 => n1558, C2 => n1157, ZN => n3796);
   U3578 : AOI221_X1 port map( B1 => n751, B2 => REGISTERS_78_25_port, C1 => 
                           n748, C2 => REGISTERS_77_25_port, A => n3805, ZN => 
                           n3799);
   U3579 : OAI222_X1 port map( A1 => n2646, A2 => n745, B1 => n2678, B2 => n742
                           , C1 => n2614, C2 => n739, ZN => n3805);
   U3580 : AOI221_X1 port map( B1 => n457, B2 => REGISTERS_45_26_port, C1 => 
                           n454, C2 => REGISTERS_44_26_port, A => n5198, ZN => 
                           n5192);
   U3581 : OAI222_X1 port map( A1 => n1589, A2 => n451, B1 => n1621, B2 => n448
                           , C1 => n1557, C2 => n445, ZN => n5198);
   U3582 : AOI221_X1 port map( B1 => n39, B2 => REGISTERS_78_26_port, C1 => n36
                           , C2 => REGISTERS_77_26_port, A => n5207, ZN => 
                           n5201);
   U3583 : OAI222_X1 port map( A1 => n2645, A2 => n33, B1 => n2677, B2 => n30, 
                           C1 => n2613, C2 => n27, ZN => n5207);
   U3584 : AOI221_X1 port map( B1 => n1169, B2 => REGISTERS_45_26_port, C1 => 
                           n1166, C2 => REGISTERS_44_26_port, A => n3755, ZN =>
                           n3749);
   U3585 : OAI222_X1 port map( A1 => n1589, A2 => n1163, B1 => n1621, B2 => 
                           n1160, C1 => n1557, C2 => n1157, ZN => n3755);
   U3586 : AOI221_X1 port map( B1 => n751, B2 => REGISTERS_78_26_port, C1 => 
                           n748, C2 => REGISTERS_77_26_port, A => n3764, ZN => 
                           n3758);
   U3587 : OAI222_X1 port map( A1 => n2645, A2 => n745, B1 => n2677, B2 => n742
                           , C1 => n2613, C2 => n739, ZN => n3764);
   U3588 : AOI221_X1 port map( B1 => n457, B2 => REGISTERS_45_27_port, C1 => 
                           n454, C2 => REGISTERS_44_27_port, A => n5157, ZN => 
                           n5151);
   U3589 : OAI222_X1 port map( A1 => n1588, A2 => n451, B1 => n1620, B2 => n448
                           , C1 => n1556, C2 => n445, ZN => n5157);
   U3590 : AOI221_X1 port map( B1 => n39, B2 => REGISTERS_78_27_port, C1 => n36
                           , C2 => REGISTERS_77_27_port, A => n5166, ZN => 
                           n5160);
   U3591 : OAI222_X1 port map( A1 => n2644, A2 => n33, B1 => n2676, B2 => n30, 
                           C1 => n2612, C2 => n27, ZN => n5166);
   U3592 : AOI221_X1 port map( B1 => n1169, B2 => REGISTERS_45_27_port, C1 => 
                           n1166, C2 => REGISTERS_44_27_port, A => n3714, ZN =>
                           n3708);
   U3593 : OAI222_X1 port map( A1 => n1588, A2 => n1163, B1 => n1620, B2 => 
                           n1160, C1 => n1556, C2 => n1157, ZN => n3714);
   U3594 : AOI221_X1 port map( B1 => n751, B2 => REGISTERS_78_27_port, C1 => 
                           n748, C2 => REGISTERS_77_27_port, A => n3723, ZN => 
                           n3717);
   U3595 : OAI222_X1 port map( A1 => n2644, A2 => n745, B1 => n2676, B2 => n742
                           , C1 => n2612, C2 => n739, ZN => n3723);
   U3596 : AOI221_X1 port map( B1 => n457, B2 => REGISTERS_45_28_port, C1 => 
                           n454, C2 => REGISTERS_44_28_port, A => n5116, ZN => 
                           n5110);
   U3597 : OAI222_X1 port map( A1 => n1587, A2 => n451, B1 => n1619, B2 => n448
                           , C1 => n1555, C2 => n445, ZN => n5116);
   U3598 : AOI221_X1 port map( B1 => n39, B2 => REGISTERS_78_28_port, C1 => n36
                           , C2 => REGISTERS_77_28_port, A => n5125, ZN => 
                           n5119);
   U3599 : OAI222_X1 port map( A1 => n2643, A2 => n33, B1 => n2675, B2 => n30, 
                           C1 => n2611, C2 => n27, ZN => n5125);
   U3600 : AOI221_X1 port map( B1 => n1169, B2 => REGISTERS_45_28_port, C1 => 
                           n1166, C2 => REGISTERS_44_28_port, A => n3673, ZN =>
                           n3667);
   U3601 : OAI222_X1 port map( A1 => n1587, A2 => n1163, B1 => n1619, B2 => 
                           n1160, C1 => n1555, C2 => n1157, ZN => n3673);
   U3602 : AOI221_X1 port map( B1 => n751, B2 => REGISTERS_78_28_port, C1 => 
                           n748, C2 => REGISTERS_77_28_port, A => n3682, ZN => 
                           n3676);
   U3603 : OAI222_X1 port map( A1 => n2643, A2 => n745, B1 => n2675, B2 => n742
                           , C1 => n2611, C2 => n739, ZN => n3682);
   U3604 : AOI221_X1 port map( B1 => n457, B2 => REGISTERS_45_29_port, C1 => 
                           n454, C2 => REGISTERS_44_29_port, A => n5075, ZN => 
                           n5069);
   U3605 : OAI222_X1 port map( A1 => n1586, A2 => n451, B1 => n1618, B2 => n448
                           , C1 => n1554, C2 => n445, ZN => n5075);
   U3606 : AOI221_X1 port map( B1 => n39, B2 => REGISTERS_78_29_port, C1 => n36
                           , C2 => REGISTERS_77_29_port, A => n5084, ZN => 
                           n5078);
   U3607 : OAI222_X1 port map( A1 => n2642, A2 => n33, B1 => n2674, B2 => n30, 
                           C1 => n2610, C2 => n27, ZN => n5084);
   U3608 : AOI221_X1 port map( B1 => n1169, B2 => REGISTERS_45_29_port, C1 => 
                           n1166, C2 => REGISTERS_44_29_port, A => n3632, ZN =>
                           n3626);
   U3609 : OAI222_X1 port map( A1 => n1586, A2 => n1163, B1 => n1618, B2 => 
                           n1160, C1 => n1554, C2 => n1157, ZN => n3632);
   U3610 : AOI221_X1 port map( B1 => n751, B2 => REGISTERS_78_29_port, C1 => 
                           n748, C2 => REGISTERS_77_29_port, A => n3641, ZN => 
                           n3635);
   U3611 : OAI222_X1 port map( A1 => n2642, A2 => n745, B1 => n2674, B2 => n742
                           , C1 => n2610, C2 => n739, ZN => n3641);
   U3612 : AOI221_X1 port map( B1 => n457, B2 => REGISTERS_45_30_port, C1 => 
                           n454, C2 => REGISTERS_44_30_port, A => n5034, ZN => 
                           n5028);
   U3613 : OAI222_X1 port map( A1 => n1585, A2 => n451, B1 => n1617, B2 => n448
                           , C1 => n1553, C2 => n445, ZN => n5034);
   U3614 : AOI221_X1 port map( B1 => n39, B2 => REGISTERS_78_30_port, C1 => n36
                           , C2 => REGISTERS_77_30_port, A => n5043, ZN => 
                           n5037);
   U3615 : OAI222_X1 port map( A1 => n2641, A2 => n33, B1 => n2673, B2 => n30, 
                           C1 => n2609, C2 => n27, ZN => n5043);
   U3616 : AOI221_X1 port map( B1 => n1169, B2 => REGISTERS_45_30_port, C1 => 
                           n1166, C2 => REGISTERS_44_30_port, A => n3591, ZN =>
                           n3585);
   U3617 : OAI222_X1 port map( A1 => n1585, A2 => n1163, B1 => n1617, B2 => 
                           n1160, C1 => n1553, C2 => n1157, ZN => n3591);
   U3618 : AOI221_X1 port map( B1 => n751, B2 => REGISTERS_78_30_port, C1 => 
                           n748, C2 => REGISTERS_77_30_port, A => n3600, ZN => 
                           n3594);
   U3619 : OAI222_X1 port map( A1 => n2641, A2 => n745, B1 => n2673, B2 => n742
                           , C1 => n2609, C2 => n739, ZN => n3600);
   U3620 : AOI221_X1 port map( B1 => n457, B2 => REGISTERS_45_31_port, C1 => 
                           n454, C2 => REGISTERS_44_31_port, A => n4962, ZN => 
                           n4943);
   U3621 : OAI222_X1 port map( A1 => n1584, A2 => n451, B1 => n1616, B2 => n448
                           , C1 => n1552, C2 => n445, ZN => n4962);
   U3622 : AOI221_X1 port map( B1 => n39, B2 => REGISTERS_78_31_port, C1 => n36
                           , C2 => REGISTERS_77_31_port, A => n4993, ZN => 
                           n4974);
   U3623 : OAI222_X1 port map( A1 => n2640, A2 => n33, B1 => n2672, B2 => n30, 
                           C1 => n2608, C2 => n27, ZN => n4993);
   U3624 : AOI221_X1 port map( B1 => n1169, B2 => REGISTERS_45_31_port, C1 => 
                           n1166, C2 => REGISTERS_44_31_port, A => n3519, ZN =>
                           n3500);
   U3625 : OAI222_X1 port map( A1 => n1584, A2 => n1163, B1 => n1616, B2 => 
                           n1160, C1 => n1552, C2 => n1157, ZN => n3519);
   U3626 : AOI221_X1 port map( B1 => n751, B2 => REGISTERS_78_31_port, C1 => 
                           n748, C2 => REGISTERS_77_31_port, A => n3550, ZN => 
                           n3531);
   U3627 : OAI222_X1 port map( A1 => n2640, A2 => n745, B1 => n2672, B2 => n742
                           , C1 => n2608, C2 => n739, ZN => n3550);
   U3628 : AND3_X1 port map( A1 => WR, A2 => ENABLE, A3 => wr_signal, ZN => 
                           n3106);
   U3629 : OAI22_X1 port map( A1 => n87, A2 => n718, B1 => n119, B2 => n715, ZN
                           => n5261);
   U3630 : OAI22_X1 port map( A1 => n791, A2 => n652, B1 => n823, B2 => n649, 
                           ZN => n5270);
   U3631 : OAI22_X1 port map( A1 => n87, A2 => n1430, B1 => n119, B2 => n1427, 
                           ZN => n3818);
   U3632 : OAI22_X1 port map( A1 => n791, A2 => n1364, B1 => n823, B2 => n1361,
                           ZN => n3827);
   U3633 : OAI22_X1 port map( A1 => n86, A2 => n718, B1 => n118, B2 => n715, ZN
                           => n5220);
   U3634 : OAI22_X1 port map( A1 => n790, A2 => n652, B1 => n822, B2 => n649, 
                           ZN => n5229);
   U3635 : OAI22_X1 port map( A1 => n86, A2 => n1430, B1 => n118, B2 => n1427, 
                           ZN => n3777);
   U3636 : OAI22_X1 port map( A1 => n790, A2 => n1364, B1 => n822, B2 => n1361,
                           ZN => n3786);
   U3637 : OAI22_X1 port map( A1 => n85, A2 => n718, B1 => n117, B2 => n715, ZN
                           => n5179);
   U3638 : OAI22_X1 port map( A1 => n789, A2 => n652, B1 => n821, B2 => n649, 
                           ZN => n5188);
   U3639 : OAI22_X1 port map( A1 => n85, A2 => n1430, B1 => n117, B2 => n1427, 
                           ZN => n3736);
   U3640 : OAI22_X1 port map( A1 => n789, A2 => n1364, B1 => n821, B2 => n1361,
                           ZN => n3745);
   U3641 : OAI22_X1 port map( A1 => n84, A2 => n718, B1 => n116, B2 => n715, ZN
                           => n5138);
   U3642 : OAI22_X1 port map( A1 => n788, A2 => n652, B1 => n820, B2 => n649, 
                           ZN => n5147);
   U3643 : OAI22_X1 port map( A1 => n84, A2 => n1430, B1 => n116, B2 => n1427, 
                           ZN => n3695);
   U3644 : OAI22_X1 port map( A1 => n788, A2 => n1364, B1 => n820, B2 => n1361,
                           ZN => n3704);
   U3645 : OAI22_X1 port map( A1 => n83, A2 => n718, B1 => n115, B2 => n715, ZN
                           => n5097);
   U3646 : OAI22_X1 port map( A1 => n787, A2 => n652, B1 => n819, B2 => n649, 
                           ZN => n5106);
   U3647 : OAI22_X1 port map( A1 => n83, A2 => n1430, B1 => n115, B2 => n1427, 
                           ZN => n3654);
   U3648 : OAI22_X1 port map( A1 => n787, A2 => n1364, B1 => n819, B2 => n1361,
                           ZN => n3663);
   U3649 : OAI22_X1 port map( A1 => n82, A2 => n718, B1 => n114, B2 => n715, ZN
                           => n5056);
   U3650 : OAI22_X1 port map( A1 => n786, A2 => n652, B1 => n818, B2 => n649, 
                           ZN => n5065);
   U3651 : OAI22_X1 port map( A1 => n82, A2 => n1430, B1 => n114, B2 => n1427, 
                           ZN => n3613);
   U3652 : OAI22_X1 port map( A1 => n786, A2 => n1364, B1 => n818, B2 => n1361,
                           ZN => n3622);
   U3653 : OAI22_X1 port map( A1 => n81, A2 => n718, B1 => n113, B2 => n715, ZN
                           => n5015);
   U3654 : OAI22_X1 port map( A1 => n785, A2 => n652, B1 => n817, B2 => n649, 
                           ZN => n5024);
   U3655 : OAI22_X1 port map( A1 => n81, A2 => n1430, B1 => n113, B2 => n1427, 
                           ZN => n3572);
   U3656 : OAI22_X1 port map( A1 => n785, A2 => n1364, B1 => n817, B2 => n1361,
                           ZN => n3581);
   U3657 : OAI22_X1 port map( A1 => n80, A2 => n718, B1 => n112, B2 => n715, ZN
                           => n4886);
   U3658 : OAI22_X1 port map( A1 => n784, A2 => n652, B1 => n816, B2 => n649, 
                           ZN => n4917);
   U3659 : OAI22_X1 port map( A1 => n80, A2 => n1430, B1 => n112, B2 => n1427, 
                           ZN => n3443);
   U3660 : OAI22_X1 port map( A1 => n784, A2 => n1364, B1 => n816, B2 => n1361,
                           ZN => n3474);
   U3661 : OAI22_X1 port map( A1 => n111, A2 => n716, B1 => n143, B2 => n713, 
                           ZN => n6245);
   U3662 : OAI22_X1 port map( A1 => n815, A2 => n650, B1 => n847, B2 => n647, 
                           ZN => n6276);
   U3663 : OAI22_X1 port map( A1 => n111, A2 => n1428, B1 => n143, B2 => n1425,
                           ZN => n4802);
   U3664 : OAI22_X1 port map( A1 => n815, A2 => n1362, B1 => n847, B2 => n1359,
                           ZN => n4833);
   U3665 : OAI22_X1 port map( A1 => n110, A2 => n716, B1 => n142, B2 => n713, 
                           ZN => n6204);
   U3666 : OAI22_X1 port map( A1 => n814, A2 => n650, B1 => n846, B2 => n647, 
                           ZN => n6213);
   U3667 : OAI22_X1 port map( A1 => n110, A2 => n1428, B1 => n142, B2 => n1425,
                           ZN => n4761);
   U3668 : OAI22_X1 port map( A1 => n814, A2 => n1362, B1 => n846, B2 => n1359,
                           ZN => n4770);
   U3669 : OAI22_X1 port map( A1 => n109, A2 => n716, B1 => n141, B2 => n713, 
                           ZN => n6163);
   U3670 : OAI22_X1 port map( A1 => n813, A2 => n650, B1 => n845, B2 => n647, 
                           ZN => n6172);
   U3671 : OAI22_X1 port map( A1 => n109, A2 => n1428, B1 => n141, B2 => n1425,
                           ZN => n4720);
   U3672 : OAI22_X1 port map( A1 => n813, A2 => n1362, B1 => n845, B2 => n1359,
                           ZN => n4729);
   U3673 : OAI22_X1 port map( A1 => n108, A2 => n716, B1 => n140, B2 => n713, 
                           ZN => n6122);
   U3674 : OAI22_X1 port map( A1 => n812, A2 => n650, B1 => n844, B2 => n647, 
                           ZN => n6131);
   U3675 : OAI22_X1 port map( A1 => n108, A2 => n1428, B1 => n140, B2 => n1425,
                           ZN => n4679);
   U3676 : OAI22_X1 port map( A1 => n812, A2 => n1362, B1 => n844, B2 => n1359,
                           ZN => n4688);
   U3677 : OAI22_X1 port map( A1 => n107, A2 => n716, B1 => n139, B2 => n713, 
                           ZN => n6081);
   U3678 : OAI22_X1 port map( A1 => n811, A2 => n650, B1 => n843, B2 => n647, 
                           ZN => n6090);
   U3679 : OAI22_X1 port map( A1 => n107, A2 => n1428, B1 => n139, B2 => n1425,
                           ZN => n4638);
   U3680 : OAI22_X1 port map( A1 => n811, A2 => n1362, B1 => n843, B2 => n1359,
                           ZN => n4647);
   U3681 : OAI22_X1 port map( A1 => n106, A2 => n716, B1 => n138, B2 => n713, 
                           ZN => n6040);
   U3682 : OAI22_X1 port map( A1 => n810, A2 => n650, B1 => n842, B2 => n647, 
                           ZN => n6049);
   U3683 : OAI22_X1 port map( A1 => n106, A2 => n1428, B1 => n138, B2 => n1425,
                           ZN => n4597);
   U3684 : OAI22_X1 port map( A1 => n810, A2 => n1362, B1 => n842, B2 => n1359,
                           ZN => n4606);
   U3685 : OAI22_X1 port map( A1 => n105, A2 => n716, B1 => n137, B2 => n713, 
                           ZN => n5999);
   U3686 : OAI22_X1 port map( A1 => n809, A2 => n650, B1 => n841, B2 => n647, 
                           ZN => n6008);
   U3687 : OAI22_X1 port map( A1 => n105, A2 => n1428, B1 => n137, B2 => n1425,
                           ZN => n4556);
   U3688 : OAI22_X1 port map( A1 => n809, A2 => n1362, B1 => n841, B2 => n1359,
                           ZN => n4565);
   U3689 : OAI22_X1 port map( A1 => n104, A2 => n716, B1 => n136, B2 => n713, 
                           ZN => n5958);
   U3690 : OAI22_X1 port map( A1 => n808, A2 => n650, B1 => n840, B2 => n647, 
                           ZN => n5967);
   U3691 : OAI22_X1 port map( A1 => n104, A2 => n1428, B1 => n136, B2 => n1425,
                           ZN => n4515);
   U3692 : OAI22_X1 port map( A1 => n808, A2 => n1362, B1 => n840, B2 => n1359,
                           ZN => n4524);
   U3693 : OAI22_X1 port map( A1 => n103, A2 => n716, B1 => n135, B2 => n713, 
                           ZN => n5917);
   U3694 : OAI22_X1 port map( A1 => n807, A2 => n650, B1 => n839, B2 => n647, 
                           ZN => n5926);
   U3695 : OAI22_X1 port map( A1 => n103, A2 => n1428, B1 => n135, B2 => n1425,
                           ZN => n4474);
   U3696 : OAI22_X1 port map( A1 => n807, A2 => n1362, B1 => n839, B2 => n1359,
                           ZN => n4483);
   U3697 : OAI22_X1 port map( A1 => n102, A2 => n716, B1 => n134, B2 => n713, 
                           ZN => n5876);
   U3698 : OAI22_X1 port map( A1 => n806, A2 => n650, B1 => n838, B2 => n647, 
                           ZN => n5885);
   U3699 : OAI22_X1 port map( A1 => n102, A2 => n1428, B1 => n134, B2 => n1425,
                           ZN => n4433);
   U3700 : OAI22_X1 port map( A1 => n806, A2 => n1362, B1 => n838, B2 => n1359,
                           ZN => n4442);
   U3701 : OAI22_X1 port map( A1 => n101, A2 => n716, B1 => n133, B2 => n713, 
                           ZN => n5835);
   U3702 : OAI22_X1 port map( A1 => n805, A2 => n650, B1 => n837, B2 => n647, 
                           ZN => n5844);
   U3703 : OAI22_X1 port map( A1 => n101, A2 => n1428, B1 => n133, B2 => n1425,
                           ZN => n4392);
   U3704 : OAI22_X1 port map( A1 => n805, A2 => n1362, B1 => n837, B2 => n1359,
                           ZN => n4401);
   U3705 : OAI22_X1 port map( A1 => n100, A2 => n716, B1 => n132, B2 => n713, 
                           ZN => n5794);
   U3706 : OAI22_X1 port map( A1 => n804, A2 => n650, B1 => n836, B2 => n647, 
                           ZN => n5803);
   U3707 : OAI22_X1 port map( A1 => n100, A2 => n1428, B1 => n132, B2 => n1425,
                           ZN => n4351);
   U3708 : OAI22_X1 port map( A1 => n804, A2 => n1362, B1 => n836, B2 => n1359,
                           ZN => n4360);
   U3709 : OAI22_X1 port map( A1 => n99, A2 => n717, B1 => n131, B2 => n714, ZN
                           => n5753);
   U3710 : OAI22_X1 port map( A1 => n803, A2 => n651, B1 => n835, B2 => n648, 
                           ZN => n5762);
   U3711 : OAI22_X1 port map( A1 => n99, A2 => n1429, B1 => n131, B2 => n1426, 
                           ZN => n4310);
   U3712 : OAI22_X1 port map( A1 => n803, A2 => n1363, B1 => n835, B2 => n1360,
                           ZN => n4319);
   U3713 : OAI22_X1 port map( A1 => n98, A2 => n717, B1 => n130, B2 => n714, ZN
                           => n5712);
   U3714 : OAI22_X1 port map( A1 => n802, A2 => n651, B1 => n834, B2 => n648, 
                           ZN => n5721);
   U3715 : OAI22_X1 port map( A1 => n98, A2 => n1429, B1 => n130, B2 => n1426, 
                           ZN => n4269);
   U3716 : OAI22_X1 port map( A1 => n802, A2 => n1363, B1 => n834, B2 => n1360,
                           ZN => n4278);
   U3717 : OAI22_X1 port map( A1 => n97, A2 => n717, B1 => n129, B2 => n714, ZN
                           => n5671);
   U3718 : OAI22_X1 port map( A1 => n801, A2 => n651, B1 => n833, B2 => n648, 
                           ZN => n5680);
   U3719 : OAI22_X1 port map( A1 => n97, A2 => n1429, B1 => n129, B2 => n1426, 
                           ZN => n4228);
   U3720 : OAI22_X1 port map( A1 => n801, A2 => n1363, B1 => n833, B2 => n1360,
                           ZN => n4237);
   U3721 : OAI22_X1 port map( A1 => n96, A2 => n717, B1 => n128, B2 => n714, ZN
                           => n5630);
   U3722 : OAI22_X1 port map( A1 => n800, A2 => n651, B1 => n832, B2 => n648, 
                           ZN => n5639);
   U3723 : OAI22_X1 port map( A1 => n96, A2 => n1429, B1 => n128, B2 => n1426, 
                           ZN => n4187);
   U3724 : OAI22_X1 port map( A1 => n800, A2 => n1363, B1 => n832, B2 => n1360,
                           ZN => n4196);
   U3725 : OAI22_X1 port map( A1 => n95, A2 => n717, B1 => n127, B2 => n714, ZN
                           => n5589);
   U3726 : OAI22_X1 port map( A1 => n799, A2 => n651, B1 => n831, B2 => n648, 
                           ZN => n5598);
   U3727 : OAI22_X1 port map( A1 => n95, A2 => n1429, B1 => n127, B2 => n1426, 
                           ZN => n4146);
   U3728 : OAI22_X1 port map( A1 => n799, A2 => n1363, B1 => n831, B2 => n1360,
                           ZN => n4155);
   U3729 : OAI22_X1 port map( A1 => n94, A2 => n717, B1 => n126, B2 => n714, ZN
                           => n5548);
   U3730 : OAI22_X1 port map( A1 => n798, A2 => n651, B1 => n830, B2 => n648, 
                           ZN => n5557);
   U3731 : OAI22_X1 port map( A1 => n94, A2 => n1429, B1 => n126, B2 => n1426, 
                           ZN => n4105);
   U3732 : OAI22_X1 port map( A1 => n798, A2 => n1363, B1 => n830, B2 => n1360,
                           ZN => n4114);
   U3733 : OAI22_X1 port map( A1 => n93, A2 => n717, B1 => n125, B2 => n714, ZN
                           => n5507);
   U3734 : OAI22_X1 port map( A1 => n797, A2 => n651, B1 => n829, B2 => n648, 
                           ZN => n5516);
   U3735 : OAI22_X1 port map( A1 => n93, A2 => n1429, B1 => n125, B2 => n1426, 
                           ZN => n4064);
   U3736 : OAI22_X1 port map( A1 => n797, A2 => n1363, B1 => n829, B2 => n1360,
                           ZN => n4073);
   U3737 : OAI22_X1 port map( A1 => n92, A2 => n717, B1 => n124, B2 => n714, ZN
                           => n5466);
   U3738 : OAI22_X1 port map( A1 => n796, A2 => n651, B1 => n828, B2 => n648, 
                           ZN => n5475);
   U3739 : OAI22_X1 port map( A1 => n92, A2 => n1429, B1 => n124, B2 => n1426, 
                           ZN => n4023);
   U3740 : OAI22_X1 port map( A1 => n796, A2 => n1363, B1 => n828, B2 => n1360,
                           ZN => n4032);
   U3741 : OAI22_X1 port map( A1 => n91, A2 => n717, B1 => n123, B2 => n714, ZN
                           => n5425);
   U3742 : OAI22_X1 port map( A1 => n795, A2 => n651, B1 => n827, B2 => n648, 
                           ZN => n5434);
   U3743 : OAI22_X1 port map( A1 => n91, A2 => n1429, B1 => n123, B2 => n1426, 
                           ZN => n3982);
   U3744 : OAI22_X1 port map( A1 => n795, A2 => n1363, B1 => n827, B2 => n1360,
                           ZN => n3991);
   U3745 : OAI22_X1 port map( A1 => n90, A2 => n717, B1 => n122, B2 => n714, ZN
                           => n5384);
   U3746 : OAI22_X1 port map( A1 => n794, A2 => n651, B1 => n826, B2 => n648, 
                           ZN => n5393);
   U3747 : OAI22_X1 port map( A1 => n90, A2 => n1429, B1 => n122, B2 => n1426, 
                           ZN => n3941);
   U3748 : OAI22_X1 port map( A1 => n794, A2 => n1363, B1 => n826, B2 => n1360,
                           ZN => n3950);
   U3749 : OAI22_X1 port map( A1 => n89, A2 => n717, B1 => n121, B2 => n714, ZN
                           => n5343);
   U3750 : OAI22_X1 port map( A1 => n793, A2 => n651, B1 => n825, B2 => n648, 
                           ZN => n5352);
   U3751 : OAI22_X1 port map( A1 => n89, A2 => n1429, B1 => n121, B2 => n1426, 
                           ZN => n3900);
   U3752 : OAI22_X1 port map( A1 => n793, A2 => n1363, B1 => n825, B2 => n1360,
                           ZN => n3909);
   U3753 : OAI22_X1 port map( A1 => n88, A2 => n717, B1 => n120, B2 => n714, ZN
                           => n5302);
   U3754 : OAI22_X1 port map( A1 => n792, A2 => n651, B1 => n824, B2 => n648, 
                           ZN => n5311);
   U3755 : OAI22_X1 port map( A1 => n88, A2 => n1429, B1 => n120, B2 => n1426, 
                           ZN => n3859);
   U3756 : OAI22_X1 port map( A1 => n792, A2 => n1363, B1 => n824, B2 => n1360,
                           ZN => n3868);
   U3757 : NAND4_X1 port map( A1 => n6238, A2 => n6239, A3 => n6240, A4 => 
                           n6241, ZN => n6237);
   U3758 : AOI221_X1 port map( B1 => n683, B2 => REGISTERS_12_0_port, C1 => 
                           n680, C2 => REGISTERS_11_0_port, A => n6258, ZN => 
                           n6240);
   U3759 : NOR4_X1 port map( A1 => n6242, A2 => n6243, A3 => n6244, A4 => n6245
                           , ZN => n6241);
   U3760 : AOI222_X1 port map( A1 => n659, A2 => REGISTERS_16_0_port, B1 => 
                           n658, B2 => REGISTERS_18_0_port, C1 => n655, C2 => 
                           REGISTERS_17_0_port, ZN => n6238);
   U3761 : NAND4_X1 port map( A1 => n4795, A2 => n4796, A3 => n4797, A4 => 
                           n4798, ZN => n4794);
   U3762 : AOI221_X1 port map( B1 => n1395, B2 => REGISTERS_12_0_port, C1 => 
                           n1392, C2 => REGISTERS_11_0_port, A => n4815, ZN => 
                           n4797);
   U3763 : NOR4_X1 port map( A1 => n4799, A2 => n4800, A3 => n4801, A4 => n4802
                           , ZN => n4798);
   U3764 : AOI222_X1 port map( A1 => n1371, A2 => REGISTERS_16_0_port, B1 => 
                           n1370, B2 => REGISTERS_18_0_port, C1 => n1367, C2 =>
                           REGISTERS_17_0_port, ZN => n4795);
   U3765 : NAND4_X1 port map( A1 => n6197, A2 => n6198, A3 => n6199, A4 => 
                           n6200, ZN => n6196);
   U3766 : AOI221_X1 port map( B1 => n683, B2 => REGISTERS_12_1_port, C1 => 
                           n680, C2 => REGISTERS_11_1_port, A => n6205, ZN => 
                           n6199);
   U3767 : NOR4_X1 port map( A1 => n6201, A2 => n6202, A3 => n6203, A4 => n6204
                           , ZN => n6200);
   U3768 : AOI222_X1 port map( A1 => n659, A2 => REGISTERS_16_1_port, B1 => 
                           n658, B2 => REGISTERS_18_1_port, C1 => n655, C2 => 
                           REGISTERS_17_1_port, ZN => n6197);
   U3769 : NAND4_X1 port map( A1 => n4754, A2 => n4755, A3 => n4756, A4 => 
                           n4757, ZN => n4753);
   U3770 : AOI221_X1 port map( B1 => n1395, B2 => REGISTERS_12_1_port, C1 => 
                           n1392, C2 => REGISTERS_11_1_port, A => n4762, ZN => 
                           n4756);
   U3771 : NOR4_X1 port map( A1 => n4758, A2 => n4759, A3 => n4760, A4 => n4761
                           , ZN => n4757);
   U3772 : AOI222_X1 port map( A1 => n1371, A2 => REGISTERS_16_1_port, B1 => 
                           n1370, B2 => REGISTERS_18_1_port, C1 => n1367, C2 =>
                           REGISTERS_17_1_port, ZN => n4754);
   U3773 : NAND4_X1 port map( A1 => n6156, A2 => n6157, A3 => n6158, A4 => 
                           n6159, ZN => n6155);
   U3774 : AOI221_X1 port map( B1 => n683, B2 => REGISTERS_12_2_port, C1 => 
                           n680, C2 => REGISTERS_11_2_port, A => n6164, ZN => 
                           n6158);
   U3775 : NOR4_X1 port map( A1 => n6160, A2 => n6161, A3 => n6162, A4 => n6163
                           , ZN => n6159);
   U3776 : AOI222_X1 port map( A1 => n659, A2 => REGISTERS_16_2_port, B1 => 
                           n658, B2 => REGISTERS_18_2_port, C1 => n655, C2 => 
                           REGISTERS_17_2_port, ZN => n6156);
   U3777 : NAND4_X1 port map( A1 => n4713, A2 => n4714, A3 => n4715, A4 => 
                           n4716, ZN => n4712);
   U3778 : AOI221_X1 port map( B1 => n1395, B2 => REGISTERS_12_2_port, C1 => 
                           n1392, C2 => REGISTERS_11_2_port, A => n4721, ZN => 
                           n4715);
   U3779 : NOR4_X1 port map( A1 => n4717, A2 => n4718, A3 => n4719, A4 => n4720
                           , ZN => n4716);
   U3780 : AOI222_X1 port map( A1 => n1371, A2 => REGISTERS_16_2_port, B1 => 
                           n1370, B2 => REGISTERS_18_2_port, C1 => n1367, C2 =>
                           REGISTERS_17_2_port, ZN => n4713);
   U3781 : NAND4_X1 port map( A1 => n6115, A2 => n6116, A3 => n6117, A4 => 
                           n6118, ZN => n6114);
   U3782 : AOI221_X1 port map( B1 => n683, B2 => REGISTERS_12_3_port, C1 => 
                           n680, C2 => REGISTERS_11_3_port, A => n6123, ZN => 
                           n6117);
   U3783 : NOR4_X1 port map( A1 => n6119, A2 => n6120, A3 => n6121, A4 => n6122
                           , ZN => n6118);
   U3784 : AOI222_X1 port map( A1 => n659, A2 => REGISTERS_16_3_port, B1 => 
                           n658, B2 => REGISTERS_18_3_port, C1 => n655, C2 => 
                           REGISTERS_17_3_port, ZN => n6115);
   U3785 : NAND4_X1 port map( A1 => n4672, A2 => n4673, A3 => n4674, A4 => 
                           n4675, ZN => n4671);
   U3786 : AOI221_X1 port map( B1 => n1395, B2 => REGISTERS_12_3_port, C1 => 
                           n1392, C2 => REGISTERS_11_3_port, A => n4680, ZN => 
                           n4674);
   U3787 : NOR4_X1 port map( A1 => n4676, A2 => n4677, A3 => n4678, A4 => n4679
                           , ZN => n4675);
   U3788 : AOI222_X1 port map( A1 => n1371, A2 => REGISTERS_16_3_port, B1 => 
                           n1370, B2 => REGISTERS_18_3_port, C1 => n1367, C2 =>
                           REGISTERS_17_3_port, ZN => n4672);
   U3789 : NAND4_X1 port map( A1 => n6074, A2 => n6075, A3 => n6076, A4 => 
                           n6077, ZN => n6073);
   U3790 : AOI221_X1 port map( B1 => n683, B2 => REGISTERS_12_4_port, C1 => 
                           n680, C2 => REGISTERS_11_4_port, A => n6082, ZN => 
                           n6076);
   U3791 : NOR4_X1 port map( A1 => n6078, A2 => n6079, A3 => n6080, A4 => n6081
                           , ZN => n6077);
   U3792 : AOI222_X1 port map( A1 => n659, A2 => REGISTERS_16_4_port, B1 => 
                           n658, B2 => REGISTERS_18_4_port, C1 => n655, C2 => 
                           REGISTERS_17_4_port, ZN => n6074);
   U3793 : NAND4_X1 port map( A1 => n4631, A2 => n4632, A3 => n4633, A4 => 
                           n4634, ZN => n4630);
   U3794 : AOI221_X1 port map( B1 => n1395, B2 => REGISTERS_12_4_port, C1 => 
                           n1392, C2 => REGISTERS_11_4_port, A => n4639, ZN => 
                           n4633);
   U3795 : NOR4_X1 port map( A1 => n4635, A2 => n4636, A3 => n4637, A4 => n4638
                           , ZN => n4634);
   U3796 : AOI222_X1 port map( A1 => n1371, A2 => REGISTERS_16_4_port, B1 => 
                           n1370, B2 => REGISTERS_18_4_port, C1 => n1367, C2 =>
                           REGISTERS_17_4_port, ZN => n4631);
   U3797 : NAND4_X1 port map( A1 => n6033, A2 => n6034, A3 => n6035, A4 => 
                           n6036, ZN => n6032);
   U3798 : AOI221_X1 port map( B1 => n683, B2 => REGISTERS_12_5_port, C1 => 
                           n680, C2 => REGISTERS_11_5_port, A => n6041, ZN => 
                           n6035);
   U3799 : NOR4_X1 port map( A1 => n6037, A2 => n6038, A3 => n6039, A4 => n6040
                           , ZN => n6036);
   U3800 : AOI222_X1 port map( A1 => n659, A2 => REGISTERS_16_5_port, B1 => 
                           n658, B2 => REGISTERS_18_5_port, C1 => n655, C2 => 
                           REGISTERS_17_5_port, ZN => n6033);
   U3801 : NAND4_X1 port map( A1 => n4590, A2 => n4591, A3 => n4592, A4 => 
                           n4593, ZN => n4589);
   U3802 : AOI221_X1 port map( B1 => n1395, B2 => REGISTERS_12_5_port, C1 => 
                           n1392, C2 => REGISTERS_11_5_port, A => n4598, ZN => 
                           n4592);
   U3803 : NOR4_X1 port map( A1 => n4594, A2 => n4595, A3 => n4596, A4 => n4597
                           , ZN => n4593);
   U3804 : AOI222_X1 port map( A1 => n1371, A2 => REGISTERS_16_5_port, B1 => 
                           n1370, B2 => REGISTERS_18_5_port, C1 => n1367, C2 =>
                           REGISTERS_17_5_port, ZN => n4590);
   U3805 : NAND4_X1 port map( A1 => n5992, A2 => n5993, A3 => n5994, A4 => 
                           n5995, ZN => n5991);
   U3806 : AOI221_X1 port map( B1 => n683, B2 => REGISTERS_12_6_port, C1 => 
                           n680, C2 => REGISTERS_11_6_port, A => n6000, ZN => 
                           n5994);
   U3807 : NOR4_X1 port map( A1 => n5996, A2 => n5997, A3 => n5998, A4 => n5999
                           , ZN => n5995);
   U3808 : AOI222_X1 port map( A1 => n659, A2 => REGISTERS_16_6_port, B1 => 
                           n658, B2 => REGISTERS_18_6_port, C1 => n655, C2 => 
                           REGISTERS_17_6_port, ZN => n5992);
   U3809 : NAND4_X1 port map( A1 => n4549, A2 => n4550, A3 => n4551, A4 => 
                           n4552, ZN => n4548);
   U3810 : AOI221_X1 port map( B1 => n1395, B2 => REGISTERS_12_6_port, C1 => 
                           n1392, C2 => REGISTERS_11_6_port, A => n4557, ZN => 
                           n4551);
   U3811 : NOR4_X1 port map( A1 => n4553, A2 => n4554, A3 => n4555, A4 => n4556
                           , ZN => n4552);
   U3812 : AOI222_X1 port map( A1 => n1371, A2 => REGISTERS_16_6_port, B1 => 
                           n1370, B2 => REGISTERS_18_6_port, C1 => n1367, C2 =>
                           REGISTERS_17_6_port, ZN => n4549);
   U3813 : NAND4_X1 port map( A1 => n5951, A2 => n5952, A3 => n5953, A4 => 
                           n5954, ZN => n5950);
   U3814 : AOI221_X1 port map( B1 => n683, B2 => REGISTERS_12_7_port, C1 => 
                           n680, C2 => REGISTERS_11_7_port, A => n5959, ZN => 
                           n5953);
   U3815 : NOR4_X1 port map( A1 => n5955, A2 => n5956, A3 => n5957, A4 => n5958
                           , ZN => n5954);
   U3816 : AOI222_X1 port map( A1 => n659, A2 => REGISTERS_16_7_port, B1 => 
                           n658, B2 => REGISTERS_18_7_port, C1 => n655, C2 => 
                           REGISTERS_17_7_port, ZN => n5951);
   U3817 : NAND4_X1 port map( A1 => n4508, A2 => n4509, A3 => n4510, A4 => 
                           n4511, ZN => n4507);
   U3818 : AOI221_X1 port map( B1 => n1395, B2 => REGISTERS_12_7_port, C1 => 
                           n1392, C2 => REGISTERS_11_7_port, A => n4516, ZN => 
                           n4510);
   U3819 : NOR4_X1 port map( A1 => n4512, A2 => n4513, A3 => n4514, A4 => n4515
                           , ZN => n4511);
   U3820 : AOI222_X1 port map( A1 => n1371, A2 => REGISTERS_16_7_port, B1 => 
                           n1370, B2 => REGISTERS_18_7_port, C1 => n1367, C2 =>
                           REGISTERS_17_7_port, ZN => n4508);
   U3821 : NAND4_X1 port map( A1 => n5910, A2 => n5911, A3 => n5912, A4 => 
                           n5913, ZN => n5909);
   U3822 : AOI221_X1 port map( B1 => n683, B2 => REGISTERS_12_8_port, C1 => 
                           n680, C2 => REGISTERS_11_8_port, A => n5918, ZN => 
                           n5912);
   U3823 : NOR4_X1 port map( A1 => n5914, A2 => n5915, A3 => n5916, A4 => n5917
                           , ZN => n5913);
   U3824 : AOI222_X1 port map( A1 => n659, A2 => REGISTERS_16_8_port, B1 => 
                           n657, B2 => REGISTERS_18_8_port, C1 => n654, C2 => 
                           REGISTERS_17_8_port, ZN => n5910);
   U3825 : NAND4_X1 port map( A1 => n4467, A2 => n4468, A3 => n4469, A4 => 
                           n4470, ZN => n4466);
   U3826 : AOI221_X1 port map( B1 => n1395, B2 => REGISTERS_12_8_port, C1 => 
                           n1392, C2 => REGISTERS_11_8_port, A => n4475, ZN => 
                           n4469);
   U3827 : NOR4_X1 port map( A1 => n4471, A2 => n4472, A3 => n4473, A4 => n4474
                           , ZN => n4470);
   U3828 : AOI222_X1 port map( A1 => n1371, A2 => REGISTERS_16_8_port, B1 => 
                           n1369, B2 => REGISTERS_18_8_port, C1 => n1366, C2 =>
                           REGISTERS_17_8_port, ZN => n4467);
   U3829 : NAND4_X1 port map( A1 => n5869, A2 => n5870, A3 => n5871, A4 => 
                           n5872, ZN => n5868);
   U3830 : AOI221_X1 port map( B1 => n683, B2 => REGISTERS_12_9_port, C1 => 
                           n680, C2 => REGISTERS_11_9_port, A => n5877, ZN => 
                           n5871);
   U3831 : NOR4_X1 port map( A1 => n5873, A2 => n5874, A3 => n5875, A4 => n5876
                           , ZN => n5872);
   U3832 : AOI222_X1 port map( A1 => n659, A2 => REGISTERS_16_9_port, B1 => 
                           n657, B2 => REGISTERS_18_9_port, C1 => n654, C2 => 
                           REGISTERS_17_9_port, ZN => n5869);
   U3833 : NAND4_X1 port map( A1 => n4426, A2 => n4427, A3 => n4428, A4 => 
                           n4429, ZN => n4425);
   U3834 : AOI221_X1 port map( B1 => n1395, B2 => REGISTERS_12_9_port, C1 => 
                           n1392, C2 => REGISTERS_11_9_port, A => n4434, ZN => 
                           n4428);
   U3835 : NOR4_X1 port map( A1 => n4430, A2 => n4431, A3 => n4432, A4 => n4433
                           , ZN => n4429);
   U3836 : AOI222_X1 port map( A1 => n1371, A2 => REGISTERS_16_9_port, B1 => 
                           n1369, B2 => REGISTERS_18_9_port, C1 => n1366, C2 =>
                           REGISTERS_17_9_port, ZN => n4426);
   U3837 : NAND4_X1 port map( A1 => n5828, A2 => n5829, A3 => n5830, A4 => 
                           n5831, ZN => n5827);
   U3838 : AOI221_X1 port map( B1 => n683, B2 => REGISTERS_12_10_port, C1 => 
                           n680, C2 => REGISTERS_11_10_port, A => n5836, ZN => 
                           n5830);
   U3839 : NOR4_X1 port map( A1 => n5832, A2 => n5833, A3 => n5834, A4 => n5835
                           , ZN => n5831);
   U3840 : AOI222_X1 port map( A1 => n659, A2 => REGISTERS_16_10_port, B1 => 
                           n657, B2 => REGISTERS_18_10_port, C1 => n654, C2 => 
                           REGISTERS_17_10_port, ZN => n5828);
   U3841 : NAND4_X1 port map( A1 => n4385, A2 => n4386, A3 => n4387, A4 => 
                           n4388, ZN => n4384);
   U3842 : AOI221_X1 port map( B1 => n1395, B2 => REGISTERS_12_10_port, C1 => 
                           n1392, C2 => REGISTERS_11_10_port, A => n4393, ZN =>
                           n4387);
   U3843 : NOR4_X1 port map( A1 => n4389, A2 => n4390, A3 => n4391, A4 => n4392
                           , ZN => n4388);
   U3844 : AOI222_X1 port map( A1 => n1371, A2 => REGISTERS_16_10_port, B1 => 
                           n1369, B2 => REGISTERS_18_10_port, C1 => n1366, C2 
                           => REGISTERS_17_10_port, ZN => n4385);
   U3845 : NAND4_X1 port map( A1 => n5787, A2 => n5788, A3 => n5789, A4 => 
                           n5790, ZN => n5786);
   U3846 : AOI221_X1 port map( B1 => n683, B2 => REGISTERS_12_11_port, C1 => 
                           n680, C2 => REGISTERS_11_11_port, A => n5795, ZN => 
                           n5789);
   U3847 : NOR4_X1 port map( A1 => n5791, A2 => n5792, A3 => n5793, A4 => n5794
                           , ZN => n5790);
   U3848 : AOI222_X1 port map( A1 => n659, A2 => REGISTERS_16_11_port, B1 => 
                           n657, B2 => REGISTERS_18_11_port, C1 => n654, C2 => 
                           REGISTERS_17_11_port, ZN => n5787);
   U3849 : NAND4_X1 port map( A1 => n4344, A2 => n4345, A3 => n4346, A4 => 
                           n4347, ZN => n4343);
   U3850 : AOI221_X1 port map( B1 => n1395, B2 => REGISTERS_12_11_port, C1 => 
                           n1392, C2 => REGISTERS_11_11_port, A => n4352, ZN =>
                           n4346);
   U3851 : NOR4_X1 port map( A1 => n4348, A2 => n4349, A3 => n4350, A4 => n4351
                           , ZN => n4347);
   U3852 : AOI222_X1 port map( A1 => n1371, A2 => REGISTERS_16_11_port, B1 => 
                           n1369, B2 => REGISTERS_18_11_port, C1 => n1366, C2 
                           => REGISTERS_17_11_port, ZN => n4344);
   U3853 : NAND4_X1 port map( A1 => n5746, A2 => n5747, A3 => n5748, A4 => 
                           n5749, ZN => n5745);
   U3854 : AOI221_X1 port map( B1 => n684, B2 => REGISTERS_12_12_port, C1 => 
                           n681, C2 => REGISTERS_11_12_port, A => n5754, ZN => 
                           n5748);
   U3855 : NOR4_X1 port map( A1 => n5750, A2 => n5751, A3 => n5752, A4 => n5753
                           , ZN => n5749);
   U3856 : AOI222_X1 port map( A1 => n660, A2 => REGISTERS_16_12_port, B1 => 
                           n657, B2 => REGISTERS_18_12_port, C1 => n654, C2 => 
                           REGISTERS_17_12_port, ZN => n5746);
   U3857 : NAND4_X1 port map( A1 => n4303, A2 => n4304, A3 => n4305, A4 => 
                           n4306, ZN => n4302);
   U3858 : AOI221_X1 port map( B1 => n1396, B2 => REGISTERS_12_12_port, C1 => 
                           n1393, C2 => REGISTERS_11_12_port, A => n4311, ZN =>
                           n4305);
   U3859 : NOR4_X1 port map( A1 => n4307, A2 => n4308, A3 => n4309, A4 => n4310
                           , ZN => n4306);
   U3860 : AOI222_X1 port map( A1 => n1372, A2 => REGISTERS_16_12_port, B1 => 
                           n1369, B2 => REGISTERS_18_12_port, C1 => n1366, C2 
                           => REGISTERS_17_12_port, ZN => n4303);
   U3861 : NAND4_X1 port map( A1 => n5705, A2 => n5706, A3 => n5707, A4 => 
                           n5708, ZN => n5704);
   U3862 : AOI221_X1 port map( B1 => n684, B2 => REGISTERS_12_13_port, C1 => 
                           n681, C2 => REGISTERS_11_13_port, A => n5713, ZN => 
                           n5707);
   U3863 : NOR4_X1 port map( A1 => n5709, A2 => n5710, A3 => n5711, A4 => n5712
                           , ZN => n5708);
   U3864 : AOI222_X1 port map( A1 => n660, A2 => REGISTERS_16_13_port, B1 => 
                           n657, B2 => REGISTERS_18_13_port, C1 => n654, C2 => 
                           REGISTERS_17_13_port, ZN => n5705);
   U3865 : NAND4_X1 port map( A1 => n4262, A2 => n4263, A3 => n4264, A4 => 
                           n4265, ZN => n4261);
   U3866 : AOI221_X1 port map( B1 => n1396, B2 => REGISTERS_12_13_port, C1 => 
                           n1393, C2 => REGISTERS_11_13_port, A => n4270, ZN =>
                           n4264);
   U3867 : NOR4_X1 port map( A1 => n4266, A2 => n4267, A3 => n4268, A4 => n4269
                           , ZN => n4265);
   U3868 : AOI222_X1 port map( A1 => n1372, A2 => REGISTERS_16_13_port, B1 => 
                           n1369, B2 => REGISTERS_18_13_port, C1 => n1366, C2 
                           => REGISTERS_17_13_port, ZN => n4262);
   U3869 : NAND4_X1 port map( A1 => n5664, A2 => n5665, A3 => n5666, A4 => 
                           n5667, ZN => n5663);
   U3870 : AOI221_X1 port map( B1 => n684, B2 => REGISTERS_12_14_port, C1 => 
                           n681, C2 => REGISTERS_11_14_port, A => n5672, ZN => 
                           n5666);
   U3871 : NOR4_X1 port map( A1 => n5668, A2 => n5669, A3 => n5670, A4 => n5671
                           , ZN => n5667);
   U3872 : AOI222_X1 port map( A1 => n660, A2 => REGISTERS_16_14_port, B1 => 
                           n657, B2 => REGISTERS_18_14_port, C1 => n654, C2 => 
                           REGISTERS_17_14_port, ZN => n5664);
   U3873 : NAND4_X1 port map( A1 => n4221, A2 => n4222, A3 => n4223, A4 => 
                           n4224, ZN => n4220);
   U3874 : AOI221_X1 port map( B1 => n1396, B2 => REGISTERS_12_14_port, C1 => 
                           n1393, C2 => REGISTERS_11_14_port, A => n4229, ZN =>
                           n4223);
   U3875 : NOR4_X1 port map( A1 => n4225, A2 => n4226, A3 => n4227, A4 => n4228
                           , ZN => n4224);
   U3876 : AOI222_X1 port map( A1 => n1372, A2 => REGISTERS_16_14_port, B1 => 
                           n1369, B2 => REGISTERS_18_14_port, C1 => n1366, C2 
                           => REGISTERS_17_14_port, ZN => n4221);
   U3877 : NAND4_X1 port map( A1 => n5623, A2 => n5624, A3 => n5625, A4 => 
                           n5626, ZN => n5622);
   U3878 : AOI221_X1 port map( B1 => n684, B2 => REGISTERS_12_15_port, C1 => 
                           n681, C2 => REGISTERS_11_15_port, A => n5631, ZN => 
                           n5625);
   U3879 : NOR4_X1 port map( A1 => n5627, A2 => n5628, A3 => n5629, A4 => n5630
                           , ZN => n5626);
   U3880 : AOI222_X1 port map( A1 => n660, A2 => REGISTERS_16_15_port, B1 => 
                           n657, B2 => REGISTERS_18_15_port, C1 => n654, C2 => 
                           REGISTERS_17_15_port, ZN => n5623);
   U3881 : NAND4_X1 port map( A1 => n4180, A2 => n4181, A3 => n4182, A4 => 
                           n4183, ZN => n4179);
   U3882 : AOI221_X1 port map( B1 => n1396, B2 => REGISTERS_12_15_port, C1 => 
                           n1393, C2 => REGISTERS_11_15_port, A => n4188, ZN =>
                           n4182);
   U3883 : NOR4_X1 port map( A1 => n4184, A2 => n4185, A3 => n4186, A4 => n4187
                           , ZN => n4183);
   U3884 : AOI222_X1 port map( A1 => n1372, A2 => REGISTERS_16_15_port, B1 => 
                           n1369, B2 => REGISTERS_18_15_port, C1 => n1366, C2 
                           => REGISTERS_17_15_port, ZN => n4180);
   U3885 : NAND4_X1 port map( A1 => n5582, A2 => n5583, A3 => n5584, A4 => 
                           n5585, ZN => n5581);
   U3886 : AOI221_X1 port map( B1 => n684, B2 => REGISTERS_12_16_port, C1 => 
                           n681, C2 => REGISTERS_11_16_port, A => n5590, ZN => 
                           n5584);
   U3887 : NOR4_X1 port map( A1 => n5586, A2 => n5587, A3 => n5588, A4 => n5589
                           , ZN => n5585);
   U3888 : AOI222_X1 port map( A1 => n660, A2 => REGISTERS_16_16_port, B1 => 
                           n657, B2 => REGISTERS_18_16_port, C1 => n654, C2 => 
                           REGISTERS_17_16_port, ZN => n5582);
   U3889 : NAND4_X1 port map( A1 => n4139, A2 => n4140, A3 => n4141, A4 => 
                           n4142, ZN => n4138);
   U3890 : AOI221_X1 port map( B1 => n1396, B2 => REGISTERS_12_16_port, C1 => 
                           n1393, C2 => REGISTERS_11_16_port, A => n4147, ZN =>
                           n4141);
   U3891 : NOR4_X1 port map( A1 => n4143, A2 => n4144, A3 => n4145, A4 => n4146
                           , ZN => n4142);
   U3892 : AOI222_X1 port map( A1 => n1372, A2 => REGISTERS_16_16_port, B1 => 
                           n1369, B2 => REGISTERS_18_16_port, C1 => n1366, C2 
                           => REGISTERS_17_16_port, ZN => n4139);
   U3893 : NAND4_X1 port map( A1 => n5541, A2 => n5542, A3 => n5543, A4 => 
                           n5544, ZN => n5540);
   U3894 : AOI221_X1 port map( B1 => n684, B2 => REGISTERS_12_17_port, C1 => 
                           n681, C2 => REGISTERS_11_17_port, A => n5549, ZN => 
                           n5543);
   U3895 : NOR4_X1 port map( A1 => n5545, A2 => n5546, A3 => n5547, A4 => n5548
                           , ZN => n5544);
   U3896 : AOI222_X1 port map( A1 => n660, A2 => REGISTERS_16_17_port, B1 => 
                           n657, B2 => REGISTERS_18_17_port, C1 => n654, C2 => 
                           REGISTERS_17_17_port, ZN => n5541);
   U3897 : NAND4_X1 port map( A1 => n4098, A2 => n4099, A3 => n4100, A4 => 
                           n4101, ZN => n4097);
   U3898 : AOI221_X1 port map( B1 => n1396, B2 => REGISTERS_12_17_port, C1 => 
                           n1393, C2 => REGISTERS_11_17_port, A => n4106, ZN =>
                           n4100);
   U3899 : NOR4_X1 port map( A1 => n4102, A2 => n4103, A3 => n4104, A4 => n4105
                           , ZN => n4101);
   U3900 : AOI222_X1 port map( A1 => n1372, A2 => REGISTERS_16_17_port, B1 => 
                           n1369, B2 => REGISTERS_18_17_port, C1 => n1366, C2 
                           => REGISTERS_17_17_port, ZN => n4098);
   U3901 : NAND4_X1 port map( A1 => n5500, A2 => n5501, A3 => n5502, A4 => 
                           n5503, ZN => n5499);
   U3902 : AOI221_X1 port map( B1 => n684, B2 => REGISTERS_12_18_port, C1 => 
                           n681, C2 => REGISTERS_11_18_port, A => n5508, ZN => 
                           n5502);
   U3903 : NOR4_X1 port map( A1 => n5504, A2 => n5505, A3 => n5506, A4 => n5507
                           , ZN => n5503);
   U3904 : AOI222_X1 port map( A1 => n660, A2 => REGISTERS_16_18_port, B1 => 
                           n657, B2 => REGISTERS_18_18_port, C1 => n654, C2 => 
                           REGISTERS_17_18_port, ZN => n5500);
   U3905 : NAND4_X1 port map( A1 => n4057, A2 => n4058, A3 => n4059, A4 => 
                           n4060, ZN => n4056);
   U3906 : AOI221_X1 port map( B1 => n1396, B2 => REGISTERS_12_18_port, C1 => 
                           n1393, C2 => REGISTERS_11_18_port, A => n4065, ZN =>
                           n4059);
   U3907 : NOR4_X1 port map( A1 => n4061, A2 => n4062, A3 => n4063, A4 => n4064
                           , ZN => n4060);
   U3908 : AOI222_X1 port map( A1 => n1372, A2 => REGISTERS_16_18_port, B1 => 
                           n1369, B2 => REGISTERS_18_18_port, C1 => n1366, C2 
                           => REGISTERS_17_18_port, ZN => n4057);
   U3909 : NAND4_X1 port map( A1 => n5459, A2 => n5460, A3 => n5461, A4 => 
                           n5462, ZN => n5458);
   U3910 : AOI221_X1 port map( B1 => n684, B2 => REGISTERS_12_19_port, C1 => 
                           n681, C2 => REGISTERS_11_19_port, A => n5467, ZN => 
                           n5461);
   U3911 : NOR4_X1 port map( A1 => n5463, A2 => n5464, A3 => n5465, A4 => n5466
                           , ZN => n5462);
   U3912 : AOI222_X1 port map( A1 => n660, A2 => REGISTERS_16_19_port, B1 => 
                           n657, B2 => REGISTERS_18_19_port, C1 => n654, C2 => 
                           REGISTERS_17_19_port, ZN => n5459);
   U3913 : NAND4_X1 port map( A1 => n4016, A2 => n4017, A3 => n4018, A4 => 
                           n4019, ZN => n4015);
   U3914 : AOI221_X1 port map( B1 => n1396, B2 => REGISTERS_12_19_port, C1 => 
                           n1393, C2 => REGISTERS_11_19_port, A => n4024, ZN =>
                           n4018);
   U3915 : NOR4_X1 port map( A1 => n4020, A2 => n4021, A3 => n4022, A4 => n4023
                           , ZN => n4019);
   U3916 : AOI222_X1 port map( A1 => n1372, A2 => REGISTERS_16_19_port, B1 => 
                           n1369, B2 => REGISTERS_18_19_port, C1 => n1366, C2 
                           => REGISTERS_17_19_port, ZN => n4016);
   U3917 : NAND4_X1 port map( A1 => n5418, A2 => n5419, A3 => n5420, A4 => 
                           n5421, ZN => n5417);
   U3918 : AOI221_X1 port map( B1 => n684, B2 => REGISTERS_12_20_port, C1 => 
                           n681, C2 => REGISTERS_11_20_port, A => n5426, ZN => 
                           n5420);
   U3919 : NOR4_X1 port map( A1 => n5422, A2 => n5423, A3 => n5424, A4 => n5425
                           , ZN => n5421);
   U3920 : AOI222_X1 port map( A1 => n660, A2 => REGISTERS_16_20_port, B1 => 
                           n656, B2 => REGISTERS_18_20_port, C1 => n653, C2 => 
                           REGISTERS_17_20_port, ZN => n5418);
   U3921 : NAND4_X1 port map( A1 => n3975, A2 => n3976, A3 => n3977, A4 => 
                           n3978, ZN => n3974);
   U3922 : AOI221_X1 port map( B1 => n1396, B2 => REGISTERS_12_20_port, C1 => 
                           n1393, C2 => REGISTERS_11_20_port, A => n3983, ZN =>
                           n3977);
   U3923 : NOR4_X1 port map( A1 => n3979, A2 => n3980, A3 => n3981, A4 => n3982
                           , ZN => n3978);
   U3924 : AOI222_X1 port map( A1 => n1372, A2 => REGISTERS_16_20_port, B1 => 
                           n1368, B2 => REGISTERS_18_20_port, C1 => n1365, C2 
                           => REGISTERS_17_20_port, ZN => n3975);
   U3925 : NAND4_X1 port map( A1 => n5377, A2 => n5378, A3 => n5379, A4 => 
                           n5380, ZN => n5376);
   U3926 : AOI221_X1 port map( B1 => n684, B2 => REGISTERS_12_21_port, C1 => 
                           n681, C2 => REGISTERS_11_21_port, A => n5385, ZN => 
                           n5379);
   U3927 : NOR4_X1 port map( A1 => n5381, A2 => n5382, A3 => n5383, A4 => n5384
                           , ZN => n5380);
   U3928 : AOI222_X1 port map( A1 => n660, A2 => REGISTERS_16_21_port, B1 => 
                           n656, B2 => REGISTERS_18_21_port, C1 => n653, C2 => 
                           REGISTERS_17_21_port, ZN => n5377);
   U3929 : NAND4_X1 port map( A1 => n3934, A2 => n3935, A3 => n3936, A4 => 
                           n3937, ZN => n3933);
   U3930 : AOI221_X1 port map( B1 => n1396, B2 => REGISTERS_12_21_port, C1 => 
                           n1393, C2 => REGISTERS_11_21_port, A => n3942, ZN =>
                           n3936);
   U3931 : NOR4_X1 port map( A1 => n3938, A2 => n3939, A3 => n3940, A4 => n3941
                           , ZN => n3937);
   U3932 : AOI222_X1 port map( A1 => n1372, A2 => REGISTERS_16_21_port, B1 => 
                           n1368, B2 => REGISTERS_18_21_port, C1 => n1365, C2 
                           => REGISTERS_17_21_port, ZN => n3934);
   U3933 : NAND4_X1 port map( A1 => n5336, A2 => n5337, A3 => n5338, A4 => 
                           n5339, ZN => n5335);
   U3934 : AOI221_X1 port map( B1 => n684, B2 => REGISTERS_12_22_port, C1 => 
                           n681, C2 => REGISTERS_11_22_port, A => n5344, ZN => 
                           n5338);
   U3935 : NOR4_X1 port map( A1 => n5340, A2 => n5341, A3 => n5342, A4 => n5343
                           , ZN => n5339);
   U3936 : AOI222_X1 port map( A1 => n660, A2 => REGISTERS_16_22_port, B1 => 
                           n656, B2 => REGISTERS_18_22_port, C1 => n653, C2 => 
                           REGISTERS_17_22_port, ZN => n5336);
   U3937 : NAND4_X1 port map( A1 => n3893, A2 => n3894, A3 => n3895, A4 => 
                           n3896, ZN => n3892);
   U3938 : AOI221_X1 port map( B1 => n1396, B2 => REGISTERS_12_22_port, C1 => 
                           n1393, C2 => REGISTERS_11_22_port, A => n3901, ZN =>
                           n3895);
   U3939 : NOR4_X1 port map( A1 => n3897, A2 => n3898, A3 => n3899, A4 => n3900
                           , ZN => n3896);
   U3940 : AOI222_X1 port map( A1 => n1372, A2 => REGISTERS_16_22_port, B1 => 
                           n1368, B2 => REGISTERS_18_22_port, C1 => n1365, C2 
                           => REGISTERS_17_22_port, ZN => n3893);
   U3941 : NAND4_X1 port map( A1 => n5295, A2 => n5296, A3 => n5297, A4 => 
                           n5298, ZN => n5294);
   U3942 : AOI221_X1 port map( B1 => n684, B2 => REGISTERS_12_23_port, C1 => 
                           n681, C2 => REGISTERS_11_23_port, A => n5303, ZN => 
                           n5297);
   U3943 : NOR4_X1 port map( A1 => n5299, A2 => n5300, A3 => n5301, A4 => n5302
                           , ZN => n5298);
   U3944 : AOI222_X1 port map( A1 => n660, A2 => REGISTERS_16_23_port, B1 => 
                           n656, B2 => REGISTERS_18_23_port, C1 => n653, C2 => 
                           REGISTERS_17_23_port, ZN => n5295);
   U3945 : NAND4_X1 port map( A1 => n3852, A2 => n3853, A3 => n3854, A4 => 
                           n3855, ZN => n3851);
   U3946 : AOI221_X1 port map( B1 => n1396, B2 => REGISTERS_12_23_port, C1 => 
                           n1393, C2 => REGISTERS_11_23_port, A => n3860, ZN =>
                           n3854);
   U3947 : NOR4_X1 port map( A1 => n3856, A2 => n3857, A3 => n3858, A4 => n3859
                           , ZN => n3855);
   U3948 : AOI222_X1 port map( A1 => n1372, A2 => REGISTERS_16_23_port, B1 => 
                           n1368, B2 => REGISTERS_18_23_port, C1 => n1365, C2 
                           => REGISTERS_17_23_port, ZN => n3852);
   U3949 : NAND4_X1 port map( A1 => n5254, A2 => n5255, A3 => n5256, A4 => 
                           n5257, ZN => n5253);
   U3950 : AOI221_X1 port map( B1 => n685, B2 => REGISTERS_12_24_port, C1 => 
                           n682, C2 => REGISTERS_11_24_port, A => n5262, ZN => 
                           n5256);
   U3951 : NOR4_X1 port map( A1 => n5258, A2 => n5259, A3 => n5260, A4 => n5261
                           , ZN => n5257);
   U3952 : AOI222_X1 port map( A1 => n661, A2 => REGISTERS_16_24_port, B1 => 
                           n656, B2 => REGISTERS_18_24_port, C1 => n653, C2 => 
                           REGISTERS_17_24_port, ZN => n5254);
   U3953 : NAND4_X1 port map( A1 => n3811, A2 => n3812, A3 => n3813, A4 => 
                           n3814, ZN => n3810);
   U3954 : AOI221_X1 port map( B1 => n1397, B2 => REGISTERS_12_24_port, C1 => 
                           n1394, C2 => REGISTERS_11_24_port, A => n3819, ZN =>
                           n3813);
   U3955 : NOR4_X1 port map( A1 => n3815, A2 => n3816, A3 => n3817, A4 => n3818
                           , ZN => n3814);
   U3956 : AOI222_X1 port map( A1 => n1373, A2 => REGISTERS_16_24_port, B1 => 
                           n1368, B2 => REGISTERS_18_24_port, C1 => n1365, C2 
                           => REGISTERS_17_24_port, ZN => n3811);
   U3957 : NAND4_X1 port map( A1 => n5213, A2 => n5214, A3 => n5215, A4 => 
                           n5216, ZN => n5212);
   U3958 : AOI221_X1 port map( B1 => n685, B2 => REGISTERS_12_25_port, C1 => 
                           n682, C2 => REGISTERS_11_25_port, A => n5221, ZN => 
                           n5215);
   U3959 : NOR4_X1 port map( A1 => n5217, A2 => n5218, A3 => n5219, A4 => n5220
                           , ZN => n5216);
   U3960 : AOI222_X1 port map( A1 => n661, A2 => REGISTERS_16_25_port, B1 => 
                           n656, B2 => REGISTERS_18_25_port, C1 => n653, C2 => 
                           REGISTERS_17_25_port, ZN => n5213);
   U3961 : NAND4_X1 port map( A1 => n3770, A2 => n3771, A3 => n3772, A4 => 
                           n3773, ZN => n3769);
   U3962 : AOI221_X1 port map( B1 => n1397, B2 => REGISTERS_12_25_port, C1 => 
                           n1394, C2 => REGISTERS_11_25_port, A => n3778, ZN =>
                           n3772);
   U3963 : NOR4_X1 port map( A1 => n3774, A2 => n3775, A3 => n3776, A4 => n3777
                           , ZN => n3773);
   U3964 : AOI222_X1 port map( A1 => n1373, A2 => REGISTERS_16_25_port, B1 => 
                           n1368, B2 => REGISTERS_18_25_port, C1 => n1365, C2 
                           => REGISTERS_17_25_port, ZN => n3770);
   U3965 : NAND4_X1 port map( A1 => n5172, A2 => n5173, A3 => n5174, A4 => 
                           n5175, ZN => n5171);
   U3966 : AOI221_X1 port map( B1 => n685, B2 => REGISTERS_12_26_port, C1 => 
                           n682, C2 => REGISTERS_11_26_port, A => n5180, ZN => 
                           n5174);
   U3967 : NOR4_X1 port map( A1 => n5176, A2 => n5177, A3 => n5178, A4 => n5179
                           , ZN => n5175);
   U3968 : AOI222_X1 port map( A1 => n661, A2 => REGISTERS_16_26_port, B1 => 
                           n656, B2 => REGISTERS_18_26_port, C1 => n653, C2 => 
                           REGISTERS_17_26_port, ZN => n5172);
   U3969 : NAND4_X1 port map( A1 => n3729, A2 => n3730, A3 => n3731, A4 => 
                           n3732, ZN => n3728);
   U3970 : AOI221_X1 port map( B1 => n1397, B2 => REGISTERS_12_26_port, C1 => 
                           n1394, C2 => REGISTERS_11_26_port, A => n3737, ZN =>
                           n3731);
   U3971 : NOR4_X1 port map( A1 => n3733, A2 => n3734, A3 => n3735, A4 => n3736
                           , ZN => n3732);
   U3972 : AOI222_X1 port map( A1 => n1373, A2 => REGISTERS_16_26_port, B1 => 
                           n1368, B2 => REGISTERS_18_26_port, C1 => n1365, C2 
                           => REGISTERS_17_26_port, ZN => n3729);
   U3973 : NAND4_X1 port map( A1 => n5131, A2 => n5132, A3 => n5133, A4 => 
                           n5134, ZN => n5130);
   U3974 : AOI221_X1 port map( B1 => n685, B2 => REGISTERS_12_27_port, C1 => 
                           n682, C2 => REGISTERS_11_27_port, A => n5139, ZN => 
                           n5133);
   U3975 : NOR4_X1 port map( A1 => n5135, A2 => n5136, A3 => n5137, A4 => n5138
                           , ZN => n5134);
   U3976 : AOI222_X1 port map( A1 => n661, A2 => REGISTERS_16_27_port, B1 => 
                           n656, B2 => REGISTERS_18_27_port, C1 => n653, C2 => 
                           REGISTERS_17_27_port, ZN => n5131);
   U3977 : NAND4_X1 port map( A1 => n3688, A2 => n3689, A3 => n3690, A4 => 
                           n3691, ZN => n3687);
   U3978 : AOI221_X1 port map( B1 => n1397, B2 => REGISTERS_12_27_port, C1 => 
                           n1394, C2 => REGISTERS_11_27_port, A => n3696, ZN =>
                           n3690);
   U3979 : NOR4_X1 port map( A1 => n3692, A2 => n3693, A3 => n3694, A4 => n3695
                           , ZN => n3691);
   U3980 : AOI222_X1 port map( A1 => n1373, A2 => REGISTERS_16_27_port, B1 => 
                           n1368, B2 => REGISTERS_18_27_port, C1 => n1365, C2 
                           => REGISTERS_17_27_port, ZN => n3688);
   U3981 : NAND4_X1 port map( A1 => n5090, A2 => n5091, A3 => n5092, A4 => 
                           n5093, ZN => n5089);
   U3982 : AOI221_X1 port map( B1 => n685, B2 => REGISTERS_12_28_port, C1 => 
                           n682, C2 => REGISTERS_11_28_port, A => n5098, ZN => 
                           n5092);
   U3983 : NOR4_X1 port map( A1 => n5094, A2 => n5095, A3 => n5096, A4 => n5097
                           , ZN => n5093);
   U3984 : AOI222_X1 port map( A1 => n661, A2 => REGISTERS_16_28_port, B1 => 
                           n656, B2 => REGISTERS_18_28_port, C1 => n653, C2 => 
                           REGISTERS_17_28_port, ZN => n5090);
   U3985 : NAND4_X1 port map( A1 => n3647, A2 => n3648, A3 => n3649, A4 => 
                           n3650, ZN => n3646);
   U3986 : AOI221_X1 port map( B1 => n1397, B2 => REGISTERS_12_28_port, C1 => 
                           n1394, C2 => REGISTERS_11_28_port, A => n3655, ZN =>
                           n3649);
   U3987 : NOR4_X1 port map( A1 => n3651, A2 => n3652, A3 => n3653, A4 => n3654
                           , ZN => n3650);
   U3988 : AOI222_X1 port map( A1 => n1373, A2 => REGISTERS_16_28_port, B1 => 
                           n1368, B2 => REGISTERS_18_28_port, C1 => n1365, C2 
                           => REGISTERS_17_28_port, ZN => n3647);
   U3989 : NAND4_X1 port map( A1 => n5049, A2 => n5050, A3 => n5051, A4 => 
                           n5052, ZN => n5048);
   U3990 : AOI221_X1 port map( B1 => n685, B2 => REGISTERS_12_29_port, C1 => 
                           n682, C2 => REGISTERS_11_29_port, A => n5057, ZN => 
                           n5051);
   U3991 : NOR4_X1 port map( A1 => n5053, A2 => n5054, A3 => n5055, A4 => n5056
                           , ZN => n5052);
   U3992 : AOI222_X1 port map( A1 => n661, A2 => REGISTERS_16_29_port, B1 => 
                           n656, B2 => REGISTERS_18_29_port, C1 => n653, C2 => 
                           REGISTERS_17_29_port, ZN => n5049);
   U3993 : NAND4_X1 port map( A1 => n3606, A2 => n3607, A3 => n3608, A4 => 
                           n3609, ZN => n3605);
   U3994 : AOI221_X1 port map( B1 => n1397, B2 => REGISTERS_12_29_port, C1 => 
                           n1394, C2 => REGISTERS_11_29_port, A => n3614, ZN =>
                           n3608);
   U3995 : NOR4_X1 port map( A1 => n3610, A2 => n3611, A3 => n3612, A4 => n3613
                           , ZN => n3609);
   U3996 : AOI222_X1 port map( A1 => n1373, A2 => REGISTERS_16_29_port, B1 => 
                           n1368, B2 => REGISTERS_18_29_port, C1 => n1365, C2 
                           => REGISTERS_17_29_port, ZN => n3606);
   U3997 : NAND4_X1 port map( A1 => n5008, A2 => n5009, A3 => n5010, A4 => 
                           n5011, ZN => n5007);
   U3998 : AOI221_X1 port map( B1 => n685, B2 => REGISTERS_12_30_port, C1 => 
                           n682, C2 => REGISTERS_11_30_port, A => n5016, ZN => 
                           n5010);
   U3999 : NOR4_X1 port map( A1 => n5012, A2 => n5013, A3 => n5014, A4 => n5015
                           , ZN => n5011);
   U4000 : AOI222_X1 port map( A1 => n661, A2 => REGISTERS_16_30_port, B1 => 
                           n656, B2 => REGISTERS_18_30_port, C1 => n653, C2 => 
                           REGISTERS_17_30_port, ZN => n5008);
   U4001 : NAND4_X1 port map( A1 => n3565, A2 => n3566, A3 => n3567, A4 => 
                           n3568, ZN => n3564);
   U4002 : AOI221_X1 port map( B1 => n1397, B2 => REGISTERS_12_30_port, C1 => 
                           n1394, C2 => REGISTERS_11_30_port, A => n3573, ZN =>
                           n3567);
   U4003 : NOR4_X1 port map( A1 => n3569, A2 => n3570, A3 => n3571, A4 => n3572
                           , ZN => n3568);
   U4004 : AOI222_X1 port map( A1 => n1373, A2 => REGISTERS_16_30_port, B1 => 
                           n1368, B2 => REGISTERS_18_30_port, C1 => n1365, C2 
                           => REGISTERS_17_30_port, ZN => n3565);
   U4005 : NAND4_X1 port map( A1 => n4879, A2 => n4880, A3 => n4881, A4 => 
                           n4882, ZN => n4878);
   U4006 : AOI221_X1 port map( B1 => n685, B2 => REGISTERS_12_31_port, C1 => 
                           n682, C2 => REGISTERS_11_31_port, A => n4900, ZN => 
                           n4881);
   U4007 : NOR4_X1 port map( A1 => n4883, A2 => n4884, A3 => n4885, A4 => n4886
                           , ZN => n4882);
   U4008 : AOI222_X1 port map( A1 => n661, A2 => REGISTERS_16_31_port, B1 => 
                           n656, B2 => REGISTERS_18_31_port, C1 => n653, C2 => 
                           REGISTERS_17_31_port, ZN => n4879);
   U4009 : NAND4_X1 port map( A1 => n3436, A2 => n3437, A3 => n3438, A4 => 
                           n3439, ZN => n3435);
   U4010 : AOI221_X1 port map( B1 => n1397, B2 => REGISTERS_12_31_port, C1 => 
                           n1394, C2 => REGISTERS_11_31_port, A => n3457, ZN =>
                           n3438);
   U4011 : NOR4_X1 port map( A1 => n3440, A2 => n3441, A3 => n3442, A4 => n3443
                           , ZN => n3439);
   U4012 : AOI222_X1 port map( A1 => n1373, A2 => REGISTERS_16_31_port, B1 => 
                           n1368, B2 => REGISTERS_18_31_port, C1 => n1365, C2 
                           => REGISTERS_17_31_port, ZN => n3436);
   U4013 : NAND4_X1 port map( A1 => n6269, A2 => n6270, A3 => n6271, A4 => 
                           n6272, ZN => n6236);
   U4014 : AOI221_X1 port map( B1 => n617, B2 => REGISTERS_34_0_port, C1 => 
                           n614, C2 => REGISTERS_33_0_port, A => n6282, ZN => 
                           n6271);
   U4015 : NOR4_X1 port map( A1 => n6273, A2 => n6274, A3 => n6275, A4 => n6276
                           , ZN => n6272);
   U4016 : AOI222_X1 port map( A1 => n593, A2 => REGISTERS_38_0_port, B1 => 
                           n592, B2 => REGISTERS_40_0_port, C1 => n493, C2 => 
                           REGISTERS_39_0_port, ZN => n6269);
   U4017 : NAND4_X1 port map( A1 => n4826, A2 => n4827, A3 => n4828, A4 => 
                           n4829, ZN => n4793);
   U4018 : AOI221_X1 port map( B1 => n1329, B2 => REGISTERS_34_0_port, C1 => 
                           n1326, C2 => REGISTERS_33_0_port, A => n4839, ZN => 
                           n4828);
   U4019 : NOR4_X1 port map( A1 => n4830, A2 => n4831, A3 => n4832, A4 => n4833
                           , ZN => n4829);
   U4020 : AOI222_X1 port map( A1 => n1305, A2 => REGISTERS_38_0_port, B1 => 
                           n1304, B2 => REGISTERS_40_0_port, C1 => n1301, C2 =>
                           REGISTERS_39_0_port, ZN => n4826);
   U4021 : NAND4_X1 port map( A1 => n6206, A2 => n6207, A3 => n6208, A4 => 
                           n6209, ZN => n6195);
   U4022 : AOI221_X1 port map( B1 => n617, B2 => REGISTERS_34_1_port, C1 => 
                           n614, C2 => REGISTERS_33_1_port, A => n6214, ZN => 
                           n6208);
   U4023 : NOR4_X1 port map( A1 => n6210, A2 => n6211, A3 => n6212, A4 => n6213
                           , ZN => n6209);
   U4024 : AOI222_X1 port map( A1 => n593, A2 => REGISTERS_38_1_port, B1 => 
                           n592, B2 => REGISTERS_40_1_port, C1 => n493, C2 => 
                           REGISTERS_39_1_port, ZN => n6206);
   U4025 : NAND4_X1 port map( A1 => n4763, A2 => n4764, A3 => n4765, A4 => 
                           n4766, ZN => n4752);
   U4026 : AOI221_X1 port map( B1 => n1329, B2 => REGISTERS_34_1_port, C1 => 
                           n1326, C2 => REGISTERS_33_1_port, A => n4771, ZN => 
                           n4765);
   U4027 : NOR4_X1 port map( A1 => n4767, A2 => n4768, A3 => n4769, A4 => n4770
                           , ZN => n4766);
   U4028 : AOI222_X1 port map( A1 => n1305, A2 => REGISTERS_38_1_port, B1 => 
                           n1304, B2 => REGISTERS_40_1_port, C1 => n1301, C2 =>
                           REGISTERS_39_1_port, ZN => n4763);
   U4029 : NAND4_X1 port map( A1 => n6165, A2 => n6166, A3 => n6167, A4 => 
                           n6168, ZN => n6154);
   U4030 : AOI221_X1 port map( B1 => n617, B2 => REGISTERS_34_2_port, C1 => 
                           n614, C2 => REGISTERS_33_2_port, A => n6173, ZN => 
                           n6167);
   U4031 : NOR4_X1 port map( A1 => n6169, A2 => n6170, A3 => n6171, A4 => n6172
                           , ZN => n6168);
   U4032 : AOI222_X1 port map( A1 => n593, A2 => REGISTERS_38_2_port, B1 => 
                           n592, B2 => REGISTERS_40_2_port, C1 => n493, C2 => 
                           REGISTERS_39_2_port, ZN => n6165);
   U4033 : NAND4_X1 port map( A1 => n4722, A2 => n4723, A3 => n4724, A4 => 
                           n4725, ZN => n4711);
   U4034 : AOI221_X1 port map( B1 => n1329, B2 => REGISTERS_34_2_port, C1 => 
                           n1326, C2 => REGISTERS_33_2_port, A => n4730, ZN => 
                           n4724);
   U4035 : NOR4_X1 port map( A1 => n4726, A2 => n4727, A3 => n4728, A4 => n4729
                           , ZN => n4725);
   U4036 : AOI222_X1 port map( A1 => n1305, A2 => REGISTERS_38_2_port, B1 => 
                           n1304, B2 => REGISTERS_40_2_port, C1 => n1301, C2 =>
                           REGISTERS_39_2_port, ZN => n4722);
   U4037 : NAND4_X1 port map( A1 => n6124, A2 => n6125, A3 => n6126, A4 => 
                           n6127, ZN => n6113);
   U4038 : AOI221_X1 port map( B1 => n617, B2 => REGISTERS_34_3_port, C1 => 
                           n614, C2 => REGISTERS_33_3_port, A => n6132, ZN => 
                           n6126);
   U4039 : NOR4_X1 port map( A1 => n6128, A2 => n6129, A3 => n6130, A4 => n6131
                           , ZN => n6127);
   U4040 : AOI222_X1 port map( A1 => n593, A2 => REGISTERS_38_3_port, B1 => 
                           n592, B2 => REGISTERS_40_3_port, C1 => n493, C2 => 
                           REGISTERS_39_3_port, ZN => n6124);
   U4041 : NAND4_X1 port map( A1 => n4681, A2 => n4682, A3 => n4683, A4 => 
                           n4684, ZN => n4670);
   U4042 : AOI221_X1 port map( B1 => n1329, B2 => REGISTERS_34_3_port, C1 => 
                           n1326, C2 => REGISTERS_33_3_port, A => n4689, ZN => 
                           n4683);
   U4043 : NOR4_X1 port map( A1 => n4685, A2 => n4686, A3 => n4687, A4 => n4688
                           , ZN => n4684);
   U4044 : AOI222_X1 port map( A1 => n1305, A2 => REGISTERS_38_3_port, B1 => 
                           n1304, B2 => REGISTERS_40_3_port, C1 => n1301, C2 =>
                           REGISTERS_39_3_port, ZN => n4681);
   U4045 : NAND4_X1 port map( A1 => n6083, A2 => n6084, A3 => n6085, A4 => 
                           n6086, ZN => n6072);
   U4046 : AOI221_X1 port map( B1 => n617, B2 => REGISTERS_34_4_port, C1 => 
                           n614, C2 => REGISTERS_33_4_port, A => n6091, ZN => 
                           n6085);
   U4047 : NOR4_X1 port map( A1 => n6087, A2 => n6088, A3 => n6089, A4 => n6090
                           , ZN => n6086);
   U4048 : AOI222_X1 port map( A1 => n593, A2 => REGISTERS_38_4_port, B1 => 
                           n592, B2 => REGISTERS_40_4_port, C1 => n493, C2 => 
                           REGISTERS_39_4_port, ZN => n6083);
   U4049 : NAND4_X1 port map( A1 => n4640, A2 => n4641, A3 => n4642, A4 => 
                           n4643, ZN => n4629);
   U4050 : AOI221_X1 port map( B1 => n1329, B2 => REGISTERS_34_4_port, C1 => 
                           n1326, C2 => REGISTERS_33_4_port, A => n4648, ZN => 
                           n4642);
   U4051 : NOR4_X1 port map( A1 => n4644, A2 => n4645, A3 => n4646, A4 => n4647
                           , ZN => n4643);
   U4052 : AOI222_X1 port map( A1 => n1305, A2 => REGISTERS_38_4_port, B1 => 
                           n1304, B2 => REGISTERS_40_4_port, C1 => n1301, C2 =>
                           REGISTERS_39_4_port, ZN => n4640);
   U4053 : NAND4_X1 port map( A1 => n6042, A2 => n6043, A3 => n6044, A4 => 
                           n6045, ZN => n6031);
   U4054 : AOI221_X1 port map( B1 => n617, B2 => REGISTERS_34_5_port, C1 => 
                           n614, C2 => REGISTERS_33_5_port, A => n6050, ZN => 
                           n6044);
   U4055 : NOR4_X1 port map( A1 => n6046, A2 => n6047, A3 => n6048, A4 => n6049
                           , ZN => n6045);
   U4056 : AOI222_X1 port map( A1 => n593, A2 => REGISTERS_38_5_port, B1 => 
                           n592, B2 => REGISTERS_40_5_port, C1 => n493, C2 => 
                           REGISTERS_39_5_port, ZN => n6042);
   U4057 : NAND4_X1 port map( A1 => n4599, A2 => n4600, A3 => n4601, A4 => 
                           n4602, ZN => n4588);
   U4058 : AOI221_X1 port map( B1 => n1329, B2 => REGISTERS_34_5_port, C1 => 
                           n1326, C2 => REGISTERS_33_5_port, A => n4607, ZN => 
                           n4601);
   U4059 : NOR4_X1 port map( A1 => n4603, A2 => n4604, A3 => n4605, A4 => n4606
                           , ZN => n4602);
   U4060 : AOI222_X1 port map( A1 => n1305, A2 => REGISTERS_38_5_port, B1 => 
                           n1304, B2 => REGISTERS_40_5_port, C1 => n1301, C2 =>
                           REGISTERS_39_5_port, ZN => n4599);
   U4061 : NAND4_X1 port map( A1 => n6001, A2 => n6002, A3 => n6003, A4 => 
                           n6004, ZN => n5990);
   U4062 : AOI221_X1 port map( B1 => n617, B2 => REGISTERS_34_6_port, C1 => 
                           n614, C2 => REGISTERS_33_6_port, A => n6009, ZN => 
                           n6003);
   U4063 : NOR4_X1 port map( A1 => n6005, A2 => n6006, A3 => n6007, A4 => n6008
                           , ZN => n6004);
   U4064 : AOI222_X1 port map( A1 => n593, A2 => REGISTERS_38_6_port, B1 => 
                           n592, B2 => REGISTERS_40_6_port, C1 => n493, C2 => 
                           REGISTERS_39_6_port, ZN => n6001);
   U4065 : NAND4_X1 port map( A1 => n4558, A2 => n4559, A3 => n4560, A4 => 
                           n4561, ZN => n4547);
   U4066 : AOI221_X1 port map( B1 => n1329, B2 => REGISTERS_34_6_port, C1 => 
                           n1326, C2 => REGISTERS_33_6_port, A => n4566, ZN => 
                           n4560);
   U4067 : NOR4_X1 port map( A1 => n4562, A2 => n4563, A3 => n4564, A4 => n4565
                           , ZN => n4561);
   U4068 : AOI222_X1 port map( A1 => n1305, A2 => REGISTERS_38_6_port, B1 => 
                           n1304, B2 => REGISTERS_40_6_port, C1 => n1301, C2 =>
                           REGISTERS_39_6_port, ZN => n4558);
   U4069 : NAND4_X1 port map( A1 => n5960, A2 => n5961, A3 => n5962, A4 => 
                           n5963, ZN => n5949);
   U4070 : AOI221_X1 port map( B1 => n617, B2 => REGISTERS_34_7_port, C1 => 
                           n614, C2 => REGISTERS_33_7_port, A => n5968, ZN => 
                           n5962);
   U4071 : NOR4_X1 port map( A1 => n5964, A2 => n5965, A3 => n5966, A4 => n5967
                           , ZN => n5963);
   U4072 : AOI222_X1 port map( A1 => n593, A2 => REGISTERS_38_7_port, B1 => 
                           n592, B2 => REGISTERS_40_7_port, C1 => n493, C2 => 
                           REGISTERS_39_7_port, ZN => n5960);
   U4073 : NAND4_X1 port map( A1 => n4517, A2 => n4518, A3 => n4519, A4 => 
                           n4520, ZN => n4506);
   U4074 : AOI221_X1 port map( B1 => n1329, B2 => REGISTERS_34_7_port, C1 => 
                           n1326, C2 => REGISTERS_33_7_port, A => n4525, ZN => 
                           n4519);
   U4075 : NOR4_X1 port map( A1 => n4521, A2 => n4522, A3 => n4523, A4 => n4524
                           , ZN => n4520);
   U4076 : AOI222_X1 port map( A1 => n1305, A2 => REGISTERS_38_7_port, B1 => 
                           n1304, B2 => REGISTERS_40_7_port, C1 => n1301, C2 =>
                           REGISTERS_39_7_port, ZN => n4517);
   U4077 : NAND4_X1 port map( A1 => n5919, A2 => n5920, A3 => n5921, A4 => 
                           n5922, ZN => n5908);
   U4078 : AOI221_X1 port map( B1 => n617, B2 => REGISTERS_34_8_port, C1 => 
                           n614, C2 => REGISTERS_33_8_port, A => n5927, ZN => 
                           n5921);
   U4079 : NOR4_X1 port map( A1 => n5923, A2 => n5924, A3 => n5925, A4 => n5926
                           , ZN => n5922);
   U4080 : AOI222_X1 port map( A1 => n593, A2 => REGISTERS_38_8_port, B1 => 
                           n495, B2 => REGISTERS_40_8_port, C1 => n492, C2 => 
                           REGISTERS_39_8_port, ZN => n5919);
   U4081 : NAND4_X1 port map( A1 => n4476, A2 => n4477, A3 => n4478, A4 => 
                           n4479, ZN => n4465);
   U4082 : AOI221_X1 port map( B1 => n1329, B2 => REGISTERS_34_8_port, C1 => 
                           n1326, C2 => REGISTERS_33_8_port, A => n4484, ZN => 
                           n4478);
   U4083 : NOR4_X1 port map( A1 => n4480, A2 => n4481, A3 => n4482, A4 => n4483
                           , ZN => n4479);
   U4084 : AOI222_X1 port map( A1 => n1305, A2 => REGISTERS_38_8_port, B1 => 
                           n1303, B2 => REGISTERS_40_8_port, C1 => n1300, C2 =>
                           REGISTERS_39_8_port, ZN => n4476);
   U4085 : NAND4_X1 port map( A1 => n5878, A2 => n5879, A3 => n5880, A4 => 
                           n5881, ZN => n5867);
   U4086 : AOI221_X1 port map( B1 => n617, B2 => REGISTERS_34_9_port, C1 => 
                           n614, C2 => REGISTERS_33_9_port, A => n5886, ZN => 
                           n5880);
   U4087 : NOR4_X1 port map( A1 => n5882, A2 => n5883, A3 => n5884, A4 => n5885
                           , ZN => n5881);
   U4088 : AOI222_X1 port map( A1 => n593, A2 => REGISTERS_38_9_port, B1 => 
                           n495, B2 => REGISTERS_40_9_port, C1 => n492, C2 => 
                           REGISTERS_39_9_port, ZN => n5878);
   U4089 : NAND4_X1 port map( A1 => n4435, A2 => n4436, A3 => n4437, A4 => 
                           n4438, ZN => n4424);
   U4090 : AOI221_X1 port map( B1 => n1329, B2 => REGISTERS_34_9_port, C1 => 
                           n1326, C2 => REGISTERS_33_9_port, A => n4443, ZN => 
                           n4437);
   U4091 : NOR4_X1 port map( A1 => n4439, A2 => n4440, A3 => n4441, A4 => n4442
                           , ZN => n4438);
   U4092 : AOI222_X1 port map( A1 => n1305, A2 => REGISTERS_38_9_port, B1 => 
                           n1303, B2 => REGISTERS_40_9_port, C1 => n1300, C2 =>
                           REGISTERS_39_9_port, ZN => n4435);
   U4093 : NAND4_X1 port map( A1 => n5837, A2 => n5838, A3 => n5839, A4 => 
                           n5840, ZN => n5826);
   U4094 : AOI221_X1 port map( B1 => n617, B2 => REGISTERS_34_10_port, C1 => 
                           n614, C2 => REGISTERS_33_10_port, A => n5845, ZN => 
                           n5839);
   U4095 : NOR4_X1 port map( A1 => n5841, A2 => n5842, A3 => n5843, A4 => n5844
                           , ZN => n5840);
   U4096 : AOI222_X1 port map( A1 => n593, A2 => REGISTERS_38_10_port, B1 => 
                           n495, B2 => REGISTERS_40_10_port, C1 => n492, C2 => 
                           REGISTERS_39_10_port, ZN => n5837);
   U4097 : NAND4_X1 port map( A1 => n4394, A2 => n4395, A3 => n4396, A4 => 
                           n4397, ZN => n4383);
   U4098 : AOI221_X1 port map( B1 => n1329, B2 => REGISTERS_34_10_port, C1 => 
                           n1326, C2 => REGISTERS_33_10_port, A => n4402, ZN =>
                           n4396);
   U4099 : NOR4_X1 port map( A1 => n4398, A2 => n4399, A3 => n4400, A4 => n4401
                           , ZN => n4397);
   U4100 : AOI222_X1 port map( A1 => n1305, A2 => REGISTERS_38_10_port, B1 => 
                           n1303, B2 => REGISTERS_40_10_port, C1 => n1300, C2 
                           => REGISTERS_39_10_port, ZN => n4394);
   U4101 : NAND4_X1 port map( A1 => n5796, A2 => n5797, A3 => n5798, A4 => 
                           n5799, ZN => n5785);
   U4102 : AOI221_X1 port map( B1 => n617, B2 => REGISTERS_34_11_port, C1 => 
                           n614, C2 => REGISTERS_33_11_port, A => n5804, ZN => 
                           n5798);
   U4103 : NOR4_X1 port map( A1 => n5800, A2 => n5801, A3 => n5802, A4 => n5803
                           , ZN => n5799);
   U4104 : AOI222_X1 port map( A1 => n593, A2 => REGISTERS_38_11_port, B1 => 
                           n495, B2 => REGISTERS_40_11_port, C1 => n492, C2 => 
                           REGISTERS_39_11_port, ZN => n5796);
   U4105 : NAND4_X1 port map( A1 => n4353, A2 => n4354, A3 => n4355, A4 => 
                           n4356, ZN => n4342);
   U4106 : AOI221_X1 port map( B1 => n1329, B2 => REGISTERS_34_11_port, C1 => 
                           n1326, C2 => REGISTERS_33_11_port, A => n4361, ZN =>
                           n4355);
   U4107 : NOR4_X1 port map( A1 => n4357, A2 => n4358, A3 => n4359, A4 => n4360
                           , ZN => n4356);
   U4108 : AOI222_X1 port map( A1 => n1305, A2 => REGISTERS_38_11_port, B1 => 
                           n1303, B2 => REGISTERS_40_11_port, C1 => n1300, C2 
                           => REGISTERS_39_11_port, ZN => n4353);
   U4109 : NAND4_X1 port map( A1 => n5755, A2 => n5756, A3 => n5757, A4 => 
                           n5758, ZN => n5744);
   U4110 : AOI221_X1 port map( B1 => n618, B2 => REGISTERS_34_12_port, C1 => 
                           n615, C2 => REGISTERS_33_12_port, A => n5763, ZN => 
                           n5757);
   U4111 : NOR4_X1 port map( A1 => n5759, A2 => n5760, A3 => n5761, A4 => n5762
                           , ZN => n5758);
   U4112 : AOI222_X1 port map( A1 => n594, A2 => REGISTERS_38_12_port, B1 => 
                           n495, B2 => REGISTERS_40_12_port, C1 => n492, C2 => 
                           REGISTERS_39_12_port, ZN => n5755);
   U4113 : NAND4_X1 port map( A1 => n4312, A2 => n4313, A3 => n4314, A4 => 
                           n4315, ZN => n4301);
   U4114 : AOI221_X1 port map( B1 => n1330, B2 => REGISTERS_34_12_port, C1 => 
                           n1327, C2 => REGISTERS_33_12_port, A => n4320, ZN =>
                           n4314);
   U4115 : NOR4_X1 port map( A1 => n4316, A2 => n4317, A3 => n4318, A4 => n4319
                           , ZN => n4315);
   U4116 : AOI222_X1 port map( A1 => n1306, A2 => REGISTERS_38_12_port, B1 => 
                           n1303, B2 => REGISTERS_40_12_port, C1 => n1300, C2 
                           => REGISTERS_39_12_port, ZN => n4312);
   U4117 : NAND4_X1 port map( A1 => n5714, A2 => n5715, A3 => n5716, A4 => 
                           n5717, ZN => n5703);
   U4118 : AOI221_X1 port map( B1 => n618, B2 => REGISTERS_34_13_port, C1 => 
                           n615, C2 => REGISTERS_33_13_port, A => n5722, ZN => 
                           n5716);
   U4119 : NOR4_X1 port map( A1 => n5718, A2 => n5719, A3 => n5720, A4 => n5721
                           , ZN => n5717);
   U4120 : AOI222_X1 port map( A1 => n594, A2 => REGISTERS_38_13_port, B1 => 
                           n495, B2 => REGISTERS_40_13_port, C1 => n492, C2 => 
                           REGISTERS_39_13_port, ZN => n5714);
   U4121 : NAND4_X1 port map( A1 => n4271, A2 => n4272, A3 => n4273, A4 => 
                           n4274, ZN => n4260);
   U4122 : AOI221_X1 port map( B1 => n1330, B2 => REGISTERS_34_13_port, C1 => 
                           n1327, C2 => REGISTERS_33_13_port, A => n4279, ZN =>
                           n4273);
   U4123 : NOR4_X1 port map( A1 => n4275, A2 => n4276, A3 => n4277, A4 => n4278
                           , ZN => n4274);
   U4124 : AOI222_X1 port map( A1 => n1306, A2 => REGISTERS_38_13_port, B1 => 
                           n1303, B2 => REGISTERS_40_13_port, C1 => n1300, C2 
                           => REGISTERS_39_13_port, ZN => n4271);
   U4125 : NAND4_X1 port map( A1 => n5673, A2 => n5674, A3 => n5675, A4 => 
                           n5676, ZN => n5662);
   U4126 : AOI221_X1 port map( B1 => n618, B2 => REGISTERS_34_14_port, C1 => 
                           n615, C2 => REGISTERS_33_14_port, A => n5681, ZN => 
                           n5675);
   U4127 : NOR4_X1 port map( A1 => n5677, A2 => n5678, A3 => n5679, A4 => n5680
                           , ZN => n5676);
   U4128 : AOI222_X1 port map( A1 => n594, A2 => REGISTERS_38_14_port, B1 => 
                           n495, B2 => REGISTERS_40_14_port, C1 => n492, C2 => 
                           REGISTERS_39_14_port, ZN => n5673);
   U4129 : NAND4_X1 port map( A1 => n4230, A2 => n4231, A3 => n4232, A4 => 
                           n4233, ZN => n4219);
   U4130 : AOI221_X1 port map( B1 => n1330, B2 => REGISTERS_34_14_port, C1 => 
                           n1327, C2 => REGISTERS_33_14_port, A => n4238, ZN =>
                           n4232);
   U4131 : NOR4_X1 port map( A1 => n4234, A2 => n4235, A3 => n4236, A4 => n4237
                           , ZN => n4233);
   U4132 : AOI222_X1 port map( A1 => n1306, A2 => REGISTERS_38_14_port, B1 => 
                           n1303, B2 => REGISTERS_40_14_port, C1 => n1300, C2 
                           => REGISTERS_39_14_port, ZN => n4230);
   U4133 : NAND4_X1 port map( A1 => n5632, A2 => n5633, A3 => n5634, A4 => 
                           n5635, ZN => n5621);
   U4134 : AOI221_X1 port map( B1 => n618, B2 => REGISTERS_34_15_port, C1 => 
                           n615, C2 => REGISTERS_33_15_port, A => n5640, ZN => 
                           n5634);
   U4135 : NOR4_X1 port map( A1 => n5636, A2 => n5637, A3 => n5638, A4 => n5639
                           , ZN => n5635);
   U4136 : AOI222_X1 port map( A1 => n594, A2 => REGISTERS_38_15_port, B1 => 
                           n495, B2 => REGISTERS_40_15_port, C1 => n492, C2 => 
                           REGISTERS_39_15_port, ZN => n5632);
   U4137 : NAND4_X1 port map( A1 => n4189, A2 => n4190, A3 => n4191, A4 => 
                           n4192, ZN => n4178);
   U4138 : AOI221_X1 port map( B1 => n1330, B2 => REGISTERS_34_15_port, C1 => 
                           n1327, C2 => REGISTERS_33_15_port, A => n4197, ZN =>
                           n4191);
   U4139 : NOR4_X1 port map( A1 => n4193, A2 => n4194, A3 => n4195, A4 => n4196
                           , ZN => n4192);
   U4140 : AOI222_X1 port map( A1 => n1306, A2 => REGISTERS_38_15_port, B1 => 
                           n1303, B2 => REGISTERS_40_15_port, C1 => n1300, C2 
                           => REGISTERS_39_15_port, ZN => n4189);
   U4141 : NAND4_X1 port map( A1 => n5591, A2 => n5592, A3 => n5593, A4 => 
                           n5594, ZN => n5580);
   U4142 : AOI221_X1 port map( B1 => n618, B2 => REGISTERS_34_16_port, C1 => 
                           n615, C2 => REGISTERS_33_16_port, A => n5599, ZN => 
                           n5593);
   U4143 : NOR4_X1 port map( A1 => n5595, A2 => n5596, A3 => n5597, A4 => n5598
                           , ZN => n5594);
   U4144 : AOI222_X1 port map( A1 => n594, A2 => REGISTERS_38_16_port, B1 => 
                           n495, B2 => REGISTERS_40_16_port, C1 => n492, C2 => 
                           REGISTERS_39_16_port, ZN => n5591);
   U4145 : NAND4_X1 port map( A1 => n4148, A2 => n4149, A3 => n4150, A4 => 
                           n4151, ZN => n4137);
   U4146 : AOI221_X1 port map( B1 => n1330, B2 => REGISTERS_34_16_port, C1 => 
                           n1327, C2 => REGISTERS_33_16_port, A => n4156, ZN =>
                           n4150);
   U4147 : NOR4_X1 port map( A1 => n4152, A2 => n4153, A3 => n4154, A4 => n4155
                           , ZN => n4151);
   U4148 : AOI222_X1 port map( A1 => n1306, A2 => REGISTERS_38_16_port, B1 => 
                           n1303, B2 => REGISTERS_40_16_port, C1 => n1300, C2 
                           => REGISTERS_39_16_port, ZN => n4148);
   U4149 : NAND4_X1 port map( A1 => n5550, A2 => n5551, A3 => n5552, A4 => 
                           n5553, ZN => n5539);
   U4150 : AOI221_X1 port map( B1 => n618, B2 => REGISTERS_34_17_port, C1 => 
                           n615, C2 => REGISTERS_33_17_port, A => n5558, ZN => 
                           n5552);
   U4151 : NOR4_X1 port map( A1 => n5554, A2 => n5555, A3 => n5556, A4 => n5557
                           , ZN => n5553);
   U4152 : AOI222_X1 port map( A1 => n594, A2 => REGISTERS_38_17_port, B1 => 
                           n495, B2 => REGISTERS_40_17_port, C1 => n492, C2 => 
                           REGISTERS_39_17_port, ZN => n5550);
   U4153 : NAND4_X1 port map( A1 => n4107, A2 => n4108, A3 => n4109, A4 => 
                           n4110, ZN => n4096);
   U4154 : AOI221_X1 port map( B1 => n1330, B2 => REGISTERS_34_17_port, C1 => 
                           n1327, C2 => REGISTERS_33_17_port, A => n4115, ZN =>
                           n4109);
   U4155 : NOR4_X1 port map( A1 => n4111, A2 => n4112, A3 => n4113, A4 => n4114
                           , ZN => n4110);
   U4156 : AOI222_X1 port map( A1 => n1306, A2 => REGISTERS_38_17_port, B1 => 
                           n1303, B2 => REGISTERS_40_17_port, C1 => n1300, C2 
                           => REGISTERS_39_17_port, ZN => n4107);
   U4157 : NAND4_X1 port map( A1 => n5509, A2 => n5510, A3 => n5511, A4 => 
                           n5512, ZN => n5498);
   U4158 : AOI221_X1 port map( B1 => n618, B2 => REGISTERS_34_18_port, C1 => 
                           n615, C2 => REGISTERS_33_18_port, A => n5517, ZN => 
                           n5511);
   U4159 : NOR4_X1 port map( A1 => n5513, A2 => n5514, A3 => n5515, A4 => n5516
                           , ZN => n5512);
   U4160 : AOI222_X1 port map( A1 => n594, A2 => REGISTERS_38_18_port, B1 => 
                           n495, B2 => REGISTERS_40_18_port, C1 => n492, C2 => 
                           REGISTERS_39_18_port, ZN => n5509);
   U4161 : NAND4_X1 port map( A1 => n4066, A2 => n4067, A3 => n4068, A4 => 
                           n4069, ZN => n4055);
   U4162 : AOI221_X1 port map( B1 => n1330, B2 => REGISTERS_34_18_port, C1 => 
                           n1327, C2 => REGISTERS_33_18_port, A => n4074, ZN =>
                           n4068);
   U4163 : NOR4_X1 port map( A1 => n4070, A2 => n4071, A3 => n4072, A4 => n4073
                           , ZN => n4069);
   U4164 : AOI222_X1 port map( A1 => n1306, A2 => REGISTERS_38_18_port, B1 => 
                           n1303, B2 => REGISTERS_40_18_port, C1 => n1300, C2 
                           => REGISTERS_39_18_port, ZN => n4066);
   U4165 : NAND4_X1 port map( A1 => n5468, A2 => n5469, A3 => n5470, A4 => 
                           n5471, ZN => n5457);
   U4166 : AOI221_X1 port map( B1 => n618, B2 => REGISTERS_34_19_port, C1 => 
                           n615, C2 => REGISTERS_33_19_port, A => n5476, ZN => 
                           n5470);
   U4167 : NOR4_X1 port map( A1 => n5472, A2 => n5473, A3 => n5474, A4 => n5475
                           , ZN => n5471);
   U4168 : AOI222_X1 port map( A1 => n594, A2 => REGISTERS_38_19_port, B1 => 
                           n495, B2 => REGISTERS_40_19_port, C1 => n492, C2 => 
                           REGISTERS_39_19_port, ZN => n5468);
   U4169 : NAND4_X1 port map( A1 => n4025, A2 => n4026, A3 => n4027, A4 => 
                           n4028, ZN => n4014);
   U4170 : AOI221_X1 port map( B1 => n1330, B2 => REGISTERS_34_19_port, C1 => 
                           n1327, C2 => REGISTERS_33_19_port, A => n4033, ZN =>
                           n4027);
   U4171 : NOR4_X1 port map( A1 => n4029, A2 => n4030, A3 => n4031, A4 => n4032
                           , ZN => n4028);
   U4172 : AOI222_X1 port map( A1 => n1306, A2 => REGISTERS_38_19_port, B1 => 
                           n1303, B2 => REGISTERS_40_19_port, C1 => n1300, C2 
                           => REGISTERS_39_19_port, ZN => n4025);
   U4173 : NAND4_X1 port map( A1 => n5427, A2 => n5428, A3 => n5429, A4 => 
                           n5430, ZN => n5416);
   U4174 : AOI221_X1 port map( B1 => n618, B2 => REGISTERS_34_20_port, C1 => 
                           n615, C2 => REGISTERS_33_20_port, A => n5435, ZN => 
                           n5429);
   U4175 : NOR4_X1 port map( A1 => n5431, A2 => n5432, A3 => n5433, A4 => n5434
                           , ZN => n5430);
   U4176 : AOI222_X1 port map( A1 => n594, A2 => REGISTERS_38_20_port, B1 => 
                           n494, B2 => REGISTERS_40_20_port, C1 => n491, C2 => 
                           REGISTERS_39_20_port, ZN => n5427);
   U4177 : NAND4_X1 port map( A1 => n3984, A2 => n3985, A3 => n3986, A4 => 
                           n3987, ZN => n3973);
   U4178 : AOI221_X1 port map( B1 => n1330, B2 => REGISTERS_34_20_port, C1 => 
                           n1327, C2 => REGISTERS_33_20_port, A => n3992, ZN =>
                           n3986);
   U4179 : NOR4_X1 port map( A1 => n3988, A2 => n3989, A3 => n3990, A4 => n3991
                           , ZN => n3987);
   U4180 : AOI222_X1 port map( A1 => n1306, A2 => REGISTERS_38_20_port, B1 => 
                           n1302, B2 => REGISTERS_40_20_port, C1 => n1299, C2 
                           => REGISTERS_39_20_port, ZN => n3984);
   U4181 : NAND4_X1 port map( A1 => n5386, A2 => n5387, A3 => n5388, A4 => 
                           n5389, ZN => n5375);
   U4182 : AOI221_X1 port map( B1 => n618, B2 => REGISTERS_34_21_port, C1 => 
                           n615, C2 => REGISTERS_33_21_port, A => n5394, ZN => 
                           n5388);
   U4183 : NOR4_X1 port map( A1 => n5390, A2 => n5391, A3 => n5392, A4 => n5393
                           , ZN => n5389);
   U4184 : AOI222_X1 port map( A1 => n594, A2 => REGISTERS_38_21_port, B1 => 
                           n494, B2 => REGISTERS_40_21_port, C1 => n491, C2 => 
                           REGISTERS_39_21_port, ZN => n5386);
   U4185 : NAND4_X1 port map( A1 => n3943, A2 => n3944, A3 => n3945, A4 => 
                           n3946, ZN => n3932);
   U4186 : AOI221_X1 port map( B1 => n1330, B2 => REGISTERS_34_21_port, C1 => 
                           n1327, C2 => REGISTERS_33_21_port, A => n3951, ZN =>
                           n3945);
   U4187 : NOR4_X1 port map( A1 => n3947, A2 => n3948, A3 => n3949, A4 => n3950
                           , ZN => n3946);
   U4188 : AOI222_X1 port map( A1 => n1306, A2 => REGISTERS_38_21_port, B1 => 
                           n1302, B2 => REGISTERS_40_21_port, C1 => n1299, C2 
                           => REGISTERS_39_21_port, ZN => n3943);
   U4189 : NAND4_X1 port map( A1 => n5345, A2 => n5346, A3 => n5347, A4 => 
                           n5348, ZN => n5334);
   U4190 : AOI221_X1 port map( B1 => n618, B2 => REGISTERS_34_22_port, C1 => 
                           n615, C2 => REGISTERS_33_22_port, A => n5353, ZN => 
                           n5347);
   U4191 : NOR4_X1 port map( A1 => n5349, A2 => n5350, A3 => n5351, A4 => n5352
                           , ZN => n5348);
   U4192 : AOI222_X1 port map( A1 => n594, A2 => REGISTERS_38_22_port, B1 => 
                           n494, B2 => REGISTERS_40_22_port, C1 => n491, C2 => 
                           REGISTERS_39_22_port, ZN => n5345);
   U4193 : NAND4_X1 port map( A1 => n3902, A2 => n3903, A3 => n3904, A4 => 
                           n3905, ZN => n3891);
   U4194 : AOI221_X1 port map( B1 => n1330, B2 => REGISTERS_34_22_port, C1 => 
                           n1327, C2 => REGISTERS_33_22_port, A => n3910, ZN =>
                           n3904);
   U4195 : NOR4_X1 port map( A1 => n3906, A2 => n3907, A3 => n3908, A4 => n3909
                           , ZN => n3905);
   U4196 : AOI222_X1 port map( A1 => n1306, A2 => REGISTERS_38_22_port, B1 => 
                           n1302, B2 => REGISTERS_40_22_port, C1 => n1299, C2 
                           => REGISTERS_39_22_port, ZN => n3902);
   U4197 : NAND4_X1 port map( A1 => n5304, A2 => n5305, A3 => n5306, A4 => 
                           n5307, ZN => n5293);
   U4198 : AOI221_X1 port map( B1 => n618, B2 => REGISTERS_34_23_port, C1 => 
                           n615, C2 => REGISTERS_33_23_port, A => n5312, ZN => 
                           n5306);
   U4199 : NOR4_X1 port map( A1 => n5308, A2 => n5309, A3 => n5310, A4 => n5311
                           , ZN => n5307);
   U4200 : AOI222_X1 port map( A1 => n594, A2 => REGISTERS_38_23_port, B1 => 
                           n494, B2 => REGISTERS_40_23_port, C1 => n491, C2 => 
                           REGISTERS_39_23_port, ZN => n5304);
   U4201 : NAND4_X1 port map( A1 => n3861, A2 => n3862, A3 => n3863, A4 => 
                           n3864, ZN => n3850);
   U4202 : AOI221_X1 port map( B1 => n1330, B2 => REGISTERS_34_23_port, C1 => 
                           n1327, C2 => REGISTERS_33_23_port, A => n3869, ZN =>
                           n3863);
   U4203 : NOR4_X1 port map( A1 => n3865, A2 => n3866, A3 => n3867, A4 => n3868
                           , ZN => n3864);
   U4204 : AOI222_X1 port map( A1 => n1306, A2 => REGISTERS_38_23_port, B1 => 
                           n1302, B2 => REGISTERS_40_23_port, C1 => n1299, C2 
                           => REGISTERS_39_23_port, ZN => n3861);
   U4205 : NAND4_X1 port map( A1 => n5263, A2 => n5264, A3 => n5265, A4 => 
                           n5266, ZN => n5252);
   U4206 : AOI221_X1 port map( B1 => n619, B2 => REGISTERS_34_24_port, C1 => 
                           n616, C2 => REGISTERS_33_24_port, A => n5271, ZN => 
                           n5265);
   U4207 : NOR4_X1 port map( A1 => n5267, A2 => n5268, A3 => n5269, A4 => n5270
                           , ZN => n5266);
   U4208 : AOI222_X1 port map( A1 => n595, A2 => REGISTERS_38_24_port, B1 => 
                           n494, B2 => REGISTERS_40_24_port, C1 => n491, C2 => 
                           REGISTERS_39_24_port, ZN => n5263);
   U4209 : NAND4_X1 port map( A1 => n3820, A2 => n3821, A3 => n3822, A4 => 
                           n3823, ZN => n3809);
   U4210 : AOI221_X1 port map( B1 => n1331, B2 => REGISTERS_34_24_port, C1 => 
                           n1328, C2 => REGISTERS_33_24_port, A => n3828, ZN =>
                           n3822);
   U4211 : NOR4_X1 port map( A1 => n3824, A2 => n3825, A3 => n3826, A4 => n3827
                           , ZN => n3823);
   U4212 : AOI222_X1 port map( A1 => n1307, A2 => REGISTERS_38_24_port, B1 => 
                           n1302, B2 => REGISTERS_40_24_port, C1 => n1299, C2 
                           => REGISTERS_39_24_port, ZN => n3820);
   U4213 : NAND4_X1 port map( A1 => n5222, A2 => n5223, A3 => n5224, A4 => 
                           n5225, ZN => n5211);
   U4214 : AOI221_X1 port map( B1 => n619, B2 => REGISTERS_34_25_port, C1 => 
                           n616, C2 => REGISTERS_33_25_port, A => n5230, ZN => 
                           n5224);
   U4215 : NOR4_X1 port map( A1 => n5226, A2 => n5227, A3 => n5228, A4 => n5229
                           , ZN => n5225);
   U4216 : AOI222_X1 port map( A1 => n595, A2 => REGISTERS_38_25_port, B1 => 
                           n494, B2 => REGISTERS_40_25_port, C1 => n491, C2 => 
                           REGISTERS_39_25_port, ZN => n5222);
   U4217 : NAND4_X1 port map( A1 => n3779, A2 => n3780, A3 => n3781, A4 => 
                           n3782, ZN => n3768);
   U4218 : AOI221_X1 port map( B1 => n1331, B2 => REGISTERS_34_25_port, C1 => 
                           n1328, C2 => REGISTERS_33_25_port, A => n3787, ZN =>
                           n3781);
   U4219 : NOR4_X1 port map( A1 => n3783, A2 => n3784, A3 => n3785, A4 => n3786
                           , ZN => n3782);
   U4220 : AOI222_X1 port map( A1 => n1307, A2 => REGISTERS_38_25_port, B1 => 
                           n1302, B2 => REGISTERS_40_25_port, C1 => n1299, C2 
                           => REGISTERS_39_25_port, ZN => n3779);
   U4221 : NAND4_X1 port map( A1 => n5181, A2 => n5182, A3 => n5183, A4 => 
                           n5184, ZN => n5170);
   U4222 : AOI221_X1 port map( B1 => n619, B2 => REGISTERS_34_26_port, C1 => 
                           n616, C2 => REGISTERS_33_26_port, A => n5189, ZN => 
                           n5183);
   U4223 : NOR4_X1 port map( A1 => n5185, A2 => n5186, A3 => n5187, A4 => n5188
                           , ZN => n5184);
   U4224 : AOI222_X1 port map( A1 => n595, A2 => REGISTERS_38_26_port, B1 => 
                           n494, B2 => REGISTERS_40_26_port, C1 => n491, C2 => 
                           REGISTERS_39_26_port, ZN => n5181);
   U4225 : NAND4_X1 port map( A1 => n3738, A2 => n3739, A3 => n3740, A4 => 
                           n3741, ZN => n3727);
   U4226 : AOI221_X1 port map( B1 => n1331, B2 => REGISTERS_34_26_port, C1 => 
                           n1328, C2 => REGISTERS_33_26_port, A => n3746, ZN =>
                           n3740);
   U4227 : NOR4_X1 port map( A1 => n3742, A2 => n3743, A3 => n3744, A4 => n3745
                           , ZN => n3741);
   U4228 : AOI222_X1 port map( A1 => n1307, A2 => REGISTERS_38_26_port, B1 => 
                           n1302, B2 => REGISTERS_40_26_port, C1 => n1299, C2 
                           => REGISTERS_39_26_port, ZN => n3738);
   U4229 : NAND4_X1 port map( A1 => n5140, A2 => n5141, A3 => n5142, A4 => 
                           n5143, ZN => n5129);
   U4230 : AOI221_X1 port map( B1 => n619, B2 => REGISTERS_34_27_port, C1 => 
                           n616, C2 => REGISTERS_33_27_port, A => n5148, ZN => 
                           n5142);
   U4231 : NOR4_X1 port map( A1 => n5144, A2 => n5145, A3 => n5146, A4 => n5147
                           , ZN => n5143);
   U4232 : AOI222_X1 port map( A1 => n595, A2 => REGISTERS_38_27_port, B1 => 
                           n494, B2 => REGISTERS_40_27_port, C1 => n491, C2 => 
                           REGISTERS_39_27_port, ZN => n5140);
   U4233 : NAND4_X1 port map( A1 => n3697, A2 => n3698, A3 => n3699, A4 => 
                           n3700, ZN => n3686);
   U4234 : AOI221_X1 port map( B1 => n1331, B2 => REGISTERS_34_27_port, C1 => 
                           n1328, C2 => REGISTERS_33_27_port, A => n3705, ZN =>
                           n3699);
   U4235 : NOR4_X1 port map( A1 => n3701, A2 => n3702, A3 => n3703, A4 => n3704
                           , ZN => n3700);
   U4236 : AOI222_X1 port map( A1 => n1307, A2 => REGISTERS_38_27_port, B1 => 
                           n1302, B2 => REGISTERS_40_27_port, C1 => n1299, C2 
                           => REGISTERS_39_27_port, ZN => n3697);
   U4237 : NAND4_X1 port map( A1 => n5099, A2 => n5100, A3 => n5101, A4 => 
                           n5102, ZN => n5088);
   U4238 : AOI221_X1 port map( B1 => n619, B2 => REGISTERS_34_28_port, C1 => 
                           n616, C2 => REGISTERS_33_28_port, A => n5107, ZN => 
                           n5101);
   U4239 : NOR4_X1 port map( A1 => n5103, A2 => n5104, A3 => n5105, A4 => n5106
                           , ZN => n5102);
   U4240 : AOI222_X1 port map( A1 => n595, A2 => REGISTERS_38_28_port, B1 => 
                           n494, B2 => REGISTERS_40_28_port, C1 => n491, C2 => 
                           REGISTERS_39_28_port, ZN => n5099);
   U4241 : NAND4_X1 port map( A1 => n3656, A2 => n3657, A3 => n3658, A4 => 
                           n3659, ZN => n3645);
   U4242 : AOI221_X1 port map( B1 => n1331, B2 => REGISTERS_34_28_port, C1 => 
                           n1328, C2 => REGISTERS_33_28_port, A => n3664, ZN =>
                           n3658);
   U4243 : NOR4_X1 port map( A1 => n3660, A2 => n3661, A3 => n3662, A4 => n3663
                           , ZN => n3659);
   U4244 : AOI222_X1 port map( A1 => n1307, A2 => REGISTERS_38_28_port, B1 => 
                           n1302, B2 => REGISTERS_40_28_port, C1 => n1299, C2 
                           => REGISTERS_39_28_port, ZN => n3656);
   U4245 : NAND4_X1 port map( A1 => n5058, A2 => n5059, A3 => n5060, A4 => 
                           n5061, ZN => n5047);
   U4246 : AOI221_X1 port map( B1 => n619, B2 => REGISTERS_34_29_port, C1 => 
                           n616, C2 => REGISTERS_33_29_port, A => n5066, ZN => 
                           n5060);
   U4247 : NOR4_X1 port map( A1 => n5062, A2 => n5063, A3 => n5064, A4 => n5065
                           , ZN => n5061);
   U4248 : AOI222_X1 port map( A1 => n595, A2 => REGISTERS_38_29_port, B1 => 
                           n494, B2 => REGISTERS_40_29_port, C1 => n491, C2 => 
                           REGISTERS_39_29_port, ZN => n5058);
   U4249 : NAND4_X1 port map( A1 => n3615, A2 => n3616, A3 => n3617, A4 => 
                           n3618, ZN => n3604);
   U4250 : AOI221_X1 port map( B1 => n1331, B2 => REGISTERS_34_29_port, C1 => 
                           n1328, C2 => REGISTERS_33_29_port, A => n3623, ZN =>
                           n3617);
   U4251 : NOR4_X1 port map( A1 => n3619, A2 => n3620, A3 => n3621, A4 => n3622
                           , ZN => n3618);
   U4252 : AOI222_X1 port map( A1 => n1307, A2 => REGISTERS_38_29_port, B1 => 
                           n1302, B2 => REGISTERS_40_29_port, C1 => n1299, C2 
                           => REGISTERS_39_29_port, ZN => n3615);
   U4253 : NAND4_X1 port map( A1 => n5017, A2 => n5018, A3 => n5019, A4 => 
                           n5020, ZN => n5006);
   U4254 : AOI221_X1 port map( B1 => n619, B2 => REGISTERS_34_30_port, C1 => 
                           n616, C2 => REGISTERS_33_30_port, A => n5025, ZN => 
                           n5019);
   U4255 : NOR4_X1 port map( A1 => n5021, A2 => n5022, A3 => n5023, A4 => n5024
                           , ZN => n5020);
   U4256 : AOI222_X1 port map( A1 => n595, A2 => REGISTERS_38_30_port, B1 => 
                           n494, B2 => REGISTERS_40_30_port, C1 => n491, C2 => 
                           REGISTERS_39_30_port, ZN => n5017);
   U4257 : NAND4_X1 port map( A1 => n3574, A2 => n3575, A3 => n3576, A4 => 
                           n3577, ZN => n3563);
   U4258 : AOI221_X1 port map( B1 => n1331, B2 => REGISTERS_34_30_port, C1 => 
                           n1328, C2 => REGISTERS_33_30_port, A => n3582, ZN =>
                           n3576);
   U4259 : NOR4_X1 port map( A1 => n3578, A2 => n3579, A3 => n3580, A4 => n3581
                           , ZN => n3577);
   U4260 : AOI222_X1 port map( A1 => n1307, A2 => REGISTERS_38_30_port, B1 => 
                           n1302, B2 => REGISTERS_40_30_port, C1 => n1299, C2 
                           => REGISTERS_39_30_port, ZN => n3574);
   U4261 : NAND4_X1 port map( A1 => n4910, A2 => n4911, A3 => n4912, A4 => 
                           n4913, ZN => n4877);
   U4262 : AOI221_X1 port map( B1 => n619, B2 => REGISTERS_34_31_port, C1 => 
                           n616, C2 => REGISTERS_33_31_port, A => n4931, ZN => 
                           n4912);
   U4263 : NOR4_X1 port map( A1 => n4914, A2 => n4915, A3 => n4916, A4 => n4917
                           , ZN => n4913);
   U4264 : AOI222_X1 port map( A1 => n595, A2 => REGISTERS_38_31_port, B1 => 
                           n494, B2 => REGISTERS_40_31_port, C1 => n491, C2 => 
                           REGISTERS_39_31_port, ZN => n4910);
   U4265 : NAND4_X1 port map( A1 => n3467, A2 => n3468, A3 => n3469, A4 => 
                           n3470, ZN => n3434);
   U4266 : AOI221_X1 port map( B1 => n1331, B2 => REGISTERS_34_31_port, C1 => 
                           n1328, C2 => REGISTERS_33_31_port, A => n3488, ZN =>
                           n3469);
   U4267 : NOR4_X1 port map( A1 => n3471, A2 => n3472, A3 => n3473, A4 => n3474
                           , ZN => n3470);
   U4268 : AOI222_X1 port map( A1 => n1307, A2 => REGISTERS_38_31_port, B1 => 
                           n1302, B2 => REGISTERS_40_31_port, C1 => n1299, C2 
                           => REGISTERS_39_31_port, ZN => n3467);
   U4269 : OR2_X1 port map( A1 => ADD_RD1(4), A2 => ADD_RD1(3), ZN => N8430);
   U4270 : OR2_X1 port map( A1 => ADD_RD2(4), A2 => ADD_RD2(3), ZN => N8574);
   U4271 : OR2_X1 port map( A1 => ADD_WR(4), A2 => ADD_WR(3), ZN => N2166);
   U4272 : OR2_X1 port map( A1 => RD1, A2 => n3333, ZN => N8702);
   U4273 : OR2_X1 port map( A1 => RD2, A2 => n3333, ZN => N8735);
   BUSout(31) <= '0';
   BUSout(30) <= '0';
   BUSout(29) <= '0';
   BUSout(28) <= '0';
   BUSout(27) <= '0';
   BUSout(26) <= '0';
   BUSout(25) <= '0';
   BUSout(24) <= '0';
   BUSout(23) <= '0';
   BUSout(22) <= '0';
   BUSout(21) <= '0';
   BUSout(20) <= '0';
   BUSout(19) <= '0';
   BUSout(18) <= '0';
   BUSout(17) <= '0';
   BUSout(16) <= '0';
   BUSout(15) <= '0';
   BUSout(14) <= '0';
   BUSout(13) <= '0';
   BUSout(12) <= '0';
   BUSout(11) <= '0';
   BUSout(10) <= '0';
   BUSout(9) <= '0';
   BUSout(8) <= '0';
   BUSout(7) <= '0';
   BUSout(6) <= '0';
   BUSout(5) <= '0';
   BUSout(4) <= '0';
   BUSout(3) <= '0';
   BUSout(2) <= '0';
   BUSout(1) <= '0';
   BUSout(0) <= '0';
   U4306 : CLKBUF_X1 port map( A => DATAIN(0), Z => n1797);
   U4307 : CLKBUF_X1 port map( A => DATAIN(0), Z => n1798);
   U4308 : CLKBUF_X1 port map( A => DATAIN(0), Z => n1799);
   U4309 : CLKBUF_X1 port map( A => DATAIN(1), Z => n1808);
   U4310 : CLKBUF_X1 port map( A => DATAIN(1), Z => n1809);
   U4311 : CLKBUF_X1 port map( A => DATAIN(1), Z => n1810);
   U4312 : CLKBUF_X1 port map( A => DATAIN(2), Z => n1819);
   U4313 : CLKBUF_X1 port map( A => DATAIN(2), Z => n1820);
   U4314 : CLKBUF_X1 port map( A => DATAIN(2), Z => n1821);
   U4315 : CLKBUF_X1 port map( A => DATAIN(3), Z => n1830);
   U4316 : CLKBUF_X1 port map( A => DATAIN(3), Z => n1831);
   U4317 : CLKBUF_X1 port map( A => DATAIN(3), Z => n1832);
   U4318 : CLKBUF_X1 port map( A => DATAIN(4), Z => n2545);
   U4319 : CLKBUF_X1 port map( A => DATAIN(4), Z => n2546);
   U4320 : CLKBUF_X1 port map( A => DATAIN(4), Z => n2547);
   U4321 : CLKBUF_X1 port map( A => DATAIN(5), Z => n2556);
   U4322 : CLKBUF_X1 port map( A => DATAIN(5), Z => n2557);
   U4323 : CLKBUF_X1 port map( A => DATAIN(5), Z => n2558);
   U4324 : CLKBUF_X1 port map( A => DATAIN(6), Z => n2567);
   U4325 : CLKBUF_X1 port map( A => DATAIN(6), Z => n2568);
   U4326 : CLKBUF_X1 port map( A => DATAIN(6), Z => n2569);
   U4327 : CLKBUF_X1 port map( A => DATAIN(7), Z => n2578);
   U4328 : CLKBUF_X1 port map( A => DATAIN(7), Z => n2579);
   U4329 : CLKBUF_X1 port map( A => DATAIN(7), Z => n2580);
   U4330 : CLKBUF_X1 port map( A => DATAIN(8), Z => n2589);
   U4331 : CLKBUF_X1 port map( A => DATAIN(8), Z => n2590);
   U4332 : CLKBUF_X1 port map( A => DATAIN(8), Z => n2591);
   U4333 : CLKBUF_X1 port map( A => DATAIN(9), Z => n2600);
   U4334 : CLKBUF_X1 port map( A => DATAIN(9), Z => n2601);
   U4335 : CLKBUF_X1 port map( A => DATAIN(9), Z => n2602);
   U4336 : CLKBUF_X1 port map( A => DATAIN(10), Z => n2707);
   U4337 : CLKBUF_X1 port map( A => DATAIN(10), Z => n2708);
   U4338 : CLKBUF_X1 port map( A => DATAIN(10), Z => n2709);
   U4339 : CLKBUF_X1 port map( A => DATAIN(11), Z => n2718);
   U4340 : CLKBUF_X1 port map( A => DATAIN(11), Z => n2719);
   U4341 : CLKBUF_X1 port map( A => DATAIN(11), Z => n2720);
   U4342 : CLKBUF_X1 port map( A => DATAIN(12), Z => n2729);
   U4343 : CLKBUF_X1 port map( A => DATAIN(12), Z => n2730);
   U4344 : CLKBUF_X1 port map( A => DATAIN(12), Z => n2731);
   U4345 : CLKBUF_X1 port map( A => DATAIN(13), Z => n2740);
   U4346 : CLKBUF_X1 port map( A => DATAIN(13), Z => n2741);
   U4347 : CLKBUF_X1 port map( A => DATAIN(13), Z => n2742);
   U4348 : CLKBUF_X1 port map( A => DATAIN(14), Z => n2751);
   U4349 : CLKBUF_X1 port map( A => DATAIN(14), Z => n2752);
   U4350 : CLKBUF_X1 port map( A => DATAIN(14), Z => n2753);
   U4351 : CLKBUF_X1 port map( A => DATAIN(15), Z => n2762);
   U4352 : CLKBUF_X1 port map( A => DATAIN(15), Z => n2763);
   U4353 : CLKBUF_X1 port map( A => DATAIN(15), Z => n2764);
   U4354 : CLKBUF_X1 port map( A => DATAIN(16), Z => n2773);
   U4355 : CLKBUF_X1 port map( A => DATAIN(16), Z => n2774);
   U4356 : CLKBUF_X1 port map( A => DATAIN(16), Z => n2775);
   U4357 : CLKBUF_X1 port map( A => DATAIN(17), Z => n2784);
   U4358 : CLKBUF_X1 port map( A => DATAIN(17), Z => n2785);
   U4359 : CLKBUF_X1 port map( A => DATAIN(17), Z => n2786);
   U4360 : CLKBUF_X1 port map( A => DATAIN(18), Z => n2795);
   U4361 : CLKBUF_X1 port map( A => DATAIN(18), Z => n2796);
   U4362 : CLKBUF_X1 port map( A => DATAIN(18), Z => n2797);
   U4363 : CLKBUF_X1 port map( A => DATAIN(19), Z => n2806);
   U4364 : CLKBUF_X1 port map( A => DATAIN(19), Z => n2807);
   U4365 : CLKBUF_X1 port map( A => DATAIN(19), Z => n2808);
   U4366 : CLKBUF_X1 port map( A => DATAIN(20), Z => n2817);
   U4367 : CLKBUF_X1 port map( A => DATAIN(20), Z => n2818);
   U4368 : CLKBUF_X1 port map( A => DATAIN(20), Z => n2819);
   U4369 : CLKBUF_X1 port map( A => DATAIN(21), Z => n2828);
   U4370 : CLKBUF_X1 port map( A => DATAIN(21), Z => n2829);
   U4371 : CLKBUF_X1 port map( A => DATAIN(21), Z => n2830);
   U4372 : CLKBUF_X1 port map( A => DATAIN(22), Z => n2839);
   U4373 : CLKBUF_X1 port map( A => DATAIN(22), Z => n2840);
   U4374 : CLKBUF_X1 port map( A => DATAIN(22), Z => n2841);
   U4375 : CLKBUF_X1 port map( A => DATAIN(23), Z => n2850);
   U4376 : CLKBUF_X1 port map( A => DATAIN(23), Z => n2851);
   U4377 : CLKBUF_X1 port map( A => DATAIN(23), Z => n2852);
   U4378 : CLKBUF_X1 port map( A => DATAIN(24), Z => n2861);
   U4379 : CLKBUF_X1 port map( A => DATAIN(24), Z => n2862);
   U4380 : CLKBUF_X1 port map( A => DATAIN(24), Z => n2863);
   U4381 : CLKBUF_X1 port map( A => DATAIN(25), Z => n2872);
   U4382 : CLKBUF_X1 port map( A => DATAIN(25), Z => n2873);
   U4383 : CLKBUF_X1 port map( A => DATAIN(25), Z => n2874);
   U4384 : CLKBUF_X1 port map( A => DATAIN(26), Z => n2883);
   U4385 : CLKBUF_X1 port map( A => DATAIN(26), Z => n2884);
   U4386 : CLKBUF_X1 port map( A => DATAIN(26), Z => n2885);
   U4387 : CLKBUF_X1 port map( A => DATAIN(27), Z => n2894);
   U4388 : CLKBUF_X1 port map( A => DATAIN(27), Z => n2895);
   U4389 : CLKBUF_X1 port map( A => DATAIN(27), Z => n2896);
   U4390 : CLKBUF_X1 port map( A => DATAIN(28), Z => n2906);
   U4391 : CLKBUF_X1 port map( A => DATAIN(28), Z => n2907);
   U4392 : CLKBUF_X1 port map( A => DATAIN(28), Z => n2908);
   U4393 : CLKBUF_X1 port map( A => DATAIN(29), Z => n2922);
   U4394 : CLKBUF_X1 port map( A => DATAIN(29), Z => n2923);
   U4395 : CLKBUF_X1 port map( A => DATAIN(29), Z => n2924);
   U4396 : CLKBUF_X1 port map( A => DATAIN(30), Z => n2933);
   U4397 : CLKBUF_X1 port map( A => DATAIN(30), Z => n2934);
   U4398 : CLKBUF_X1 port map( A => DATAIN(30), Z => n2935);
   U4399 : CLKBUF_X1 port map( A => DATAIN(31), Z => n2944);
   U4400 : CLKBUF_X1 port map( A => DATAIN(31), Z => n2945);
   U4401 : CLKBUF_X1 port map( A => DATAIN(31), Z => n2946);
   U4402 : INV_X1 port map( A => n3302, ZN => n2956);
   U4403 : INV_X1 port map( A => n3301, ZN => n2957);
   U4404 : INV_X1 port map( A => n3301, ZN => n2958);
   U4405 : INV_X1 port map( A => n3301, ZN => n2959);
   U4406 : INV_X1 port map( A => n3301, ZN => n2960);
   U4407 : INV_X1 port map( A => n3301, ZN => n2961);
   U4408 : INV_X1 port map( A => n3301, ZN => n2962);
   U4409 : INV_X1 port map( A => n3301, ZN => n2963);
   U4410 : INV_X1 port map( A => n3300, ZN => n2964);
   U4411 : INV_X1 port map( A => n3300, ZN => n2965);
   U4412 : INV_X1 port map( A => n3300, ZN => n2966);
   U4413 : INV_X1 port map( A => n3300, ZN => n2967);
   U4414 : INV_X1 port map( A => n3300, ZN => n2968);
   U4415 : INV_X1 port map( A => n3300, ZN => n2969);
   U4416 : INV_X1 port map( A => n3300, ZN => n2970);
   U4417 : INV_X1 port map( A => n3298, ZN => n2971);
   U4418 : INV_X1 port map( A => n3298, ZN => n2972);
   U4419 : INV_X1 port map( A => n3298, ZN => n2973);
   U4420 : INV_X1 port map( A => n3298, ZN => n2974);
   U4421 : INV_X1 port map( A => n3298, ZN => n2975);
   U4422 : INV_X1 port map( A => n3298, ZN => n2976);
   U4423 : INV_X1 port map( A => n3298, ZN => n2977);
   U4424 : INV_X1 port map( A => n3297, ZN => n2978);
   U4425 : INV_X1 port map( A => n3297, ZN => n2979);
   U4426 : INV_X1 port map( A => n3297, ZN => n2980);
   U4427 : INV_X1 port map( A => n3297, ZN => n2981);
   U4428 : INV_X1 port map( A => n3297, ZN => n2982);
   U4429 : INV_X1 port map( A => n3297, ZN => n2983);
   U4430 : INV_X1 port map( A => n3297, ZN => n2984);
   U4431 : INV_X1 port map( A => n3296, ZN => n2985);
   U4432 : INV_X1 port map( A => n3296, ZN => n2986);
   U4433 : INV_X1 port map( A => n3296, ZN => n2987);
   U4434 : INV_X1 port map( A => n3296, ZN => n2988);
   U4435 : INV_X1 port map( A => n3296, ZN => n2989);
   U4436 : INV_X1 port map( A => n3296, ZN => n2990);
   U4437 : INV_X1 port map( A => n3296, ZN => n2991);
   U4438 : INV_X1 port map( A => n3294, ZN => n2992);
   U4439 : INV_X1 port map( A => n3294, ZN => n2993);
   U4440 : INV_X1 port map( A => n3294, ZN => n2994);
   U4441 : INV_X1 port map( A => n3294, ZN => n2995);
   U4442 : INV_X1 port map( A => n3294, ZN => n2997);
   U4443 : INV_X1 port map( A => n3294, ZN => n2998);
   U4444 : INV_X1 port map( A => n3293, ZN => n2999);
   U4445 : INV_X1 port map( A => n3293, ZN => n3000);
   U4446 : INV_X1 port map( A => n3293, ZN => n3001);
   U4447 : INV_X1 port map( A => n3293, ZN => n3002);
   U4448 : INV_X1 port map( A => n3293, ZN => n3003);
   U4449 : INV_X1 port map( A => n3293, ZN => n3004);
   U4450 : INV_X1 port map( A => n3293, ZN => n3005);
   U4451 : INV_X1 port map( A => n3292, ZN => n3006);
   U4452 : INV_X1 port map( A => n3292, ZN => n3007);
   U4453 : INV_X1 port map( A => n3292, ZN => n3008);
   U4454 : INV_X1 port map( A => n3292, ZN => n3009);
   U4455 : INV_X1 port map( A => n3292, ZN => n3010);
   U4456 : INV_X1 port map( A => n3292, ZN => n3011);
   U4457 : INV_X1 port map( A => n3292, ZN => n3012);
   U4458 : INV_X1 port map( A => n3290, ZN => n3013);
   U4459 : INV_X1 port map( A => n3290, ZN => n3014);
   U4460 : INV_X1 port map( A => n3290, ZN => n3015);
   U4461 : INV_X1 port map( A => n3290, ZN => n3016);
   U4462 : INV_X1 port map( A => n3290, ZN => n3017);
   U4463 : INV_X1 port map( A => n3290, ZN => n3018);
   U4464 : INV_X1 port map( A => n3290, ZN => n3019);
   U4465 : INV_X1 port map( A => n3289, ZN => n3020);
   U4466 : INV_X1 port map( A => n3289, ZN => n3021);
   U4467 : INV_X1 port map( A => n3289, ZN => n3022);
   U4468 : INV_X1 port map( A => n3289, ZN => n3023);
   U4469 : INV_X1 port map( A => n3289, ZN => n3024);
   U4470 : INV_X1 port map( A => n3289, ZN => n3025);
   U4471 : INV_X1 port map( A => n3288, ZN => n3026);
   U4472 : INV_X1 port map( A => n3288, ZN => n3027);
   U4473 : INV_X1 port map( A => n3288, ZN => n3028);
   U4474 : INV_X1 port map( A => n3288, ZN => n3031);
   U4475 : INV_X1 port map( A => n3288, ZN => n3032);
   U4476 : INV_X1 port map( A => n3288, ZN => n3034);
   U4477 : INV_X1 port map( A => n3288, ZN => n3036);
   U4478 : INV_X1 port map( A => n3286, ZN => n3037);
   U4479 : INV_X1 port map( A => n3286, ZN => n3039);
   U4480 : INV_X1 port map( A => n3286, ZN => n3041);
   U4481 : INV_X1 port map( A => n3286, ZN => n3042);
   U4482 : INV_X1 port map( A => n3286, ZN => n3044);
   U4483 : INV_X1 port map( A => n3286, ZN => n3046);
   U4484 : INV_X1 port map( A => n3294, ZN => n3047);
   U4485 : INV_X1 port map( A => n3331, ZN => n3049);
   U4486 : INV_X1 port map( A => n3331, ZN => n3051);
   U4487 : INV_X1 port map( A => n3331, ZN => n3052);
   U4488 : INV_X1 port map( A => n3331, ZN => n3054);
   U4489 : INV_X1 port map( A => n3331, ZN => n3056);
   U4490 : INV_X1 port map( A => n3331, ZN => n3057);
   U4491 : INV_X1 port map( A => n3330, ZN => n3059);
   U4492 : INV_X1 port map( A => n3331, ZN => n3061);
   U4493 : INV_X1 port map( A => n3330, ZN => n3062);
   U4494 : INV_X1 port map( A => n3330, ZN => n3064);
   U4495 : INV_X1 port map( A => n3330, ZN => n3066);
   U4496 : INV_X1 port map( A => n3330, ZN => n3067);
   U4497 : INV_X1 port map( A => n3330, ZN => n3069);
   U4498 : INV_X1 port map( A => n3330, ZN => n3071);
   U4499 : INV_X1 port map( A => n3329, ZN => n3072);
   U4500 : INV_X1 port map( A => n3329, ZN => n3074);
   U4501 : INV_X1 port map( A => n3329, ZN => n3076);
   U4502 : INV_X1 port map( A => n3329, ZN => n3077);
   U4503 : INV_X1 port map( A => n3329, ZN => n3079);
   U4504 : INV_X1 port map( A => n3329, ZN => n3081);
   U4505 : INV_X1 port map( A => n3327, ZN => n3082);
   U4506 : INV_X1 port map( A => n3329, ZN => n3084);
   U4507 : INV_X1 port map( A => n3327, ZN => n3086);
   U4508 : INV_X1 port map( A => n3327, ZN => n3087);
   U4509 : INV_X1 port map( A => n3327, ZN => n3089);
   U4510 : INV_X1 port map( A => n3327, ZN => n3091);
   U4511 : INV_X1 port map( A => n3327, ZN => n3092);
   U4512 : INV_X1 port map( A => n3327, ZN => n3094);
   U4513 : INV_X1 port map( A => n3326, ZN => n3096);
   U4514 : INV_X1 port map( A => n3326, ZN => n3097);
   U4515 : INV_X1 port map( A => n3326, ZN => n3099);
   U4516 : INV_X1 port map( A => n3326, ZN => n3101);
   U4517 : INV_X1 port map( A => n3326, ZN => n3102);
   U4518 : INV_X1 port map( A => n3326, ZN => n3104);
   U4519 : INV_X1 port map( A => n3326, ZN => n3110);
   U4520 : INV_X1 port map( A => n3325, ZN => n3111);
   U4521 : INV_X1 port map( A => n3325, ZN => n3113);
   U4522 : INV_X1 port map( A => n3325, ZN => n3115);
   U4523 : INV_X1 port map( A => n3325, ZN => n3116);
   U4524 : INV_X1 port map( A => n3325, ZN => n3118);
   U4525 : INV_X1 port map( A => n3325, ZN => n3119);
   U4526 : INV_X1 port map( A => n3325, ZN => n3120);
   U4527 : INV_X1 port map( A => n3323, ZN => n3122);
   U4528 : INV_X1 port map( A => n3323, ZN => n3123);
   U4529 : INV_X1 port map( A => n3323, ZN => n3124);
   U4530 : INV_X1 port map( A => n3323, ZN => n3126);
   U4531 : INV_X1 port map( A => n3323, ZN => n3127);
   U4532 : INV_X1 port map( A => n3323, ZN => n3128);
   U4533 : INV_X1 port map( A => n3323, ZN => n3130);
   U4534 : INV_X1 port map( A => n3322, ZN => n3131);
   U4535 : INV_X1 port map( A => n3322, ZN => n3132);
   U4536 : INV_X1 port map( A => n3322, ZN => n3134);
   U4537 : INV_X1 port map( A => n3322, ZN => n3135);
   U4538 : INV_X1 port map( A => n3322, ZN => n3136);
   U4539 : INV_X1 port map( A => n3322, ZN => n3138);
   U4540 : INV_X1 port map( A => n3322, ZN => n3139);
   U4541 : INV_X1 port map( A => n3321, ZN => n3140);
   U4542 : INV_X1 port map( A => n3321, ZN => n3142);
   U4543 : INV_X1 port map( A => n3321, ZN => n3143);
   U4544 : INV_X1 port map( A => n3321, ZN => n3144);
   U4545 : INV_X1 port map( A => n3321, ZN => n3146);
   U4546 : INV_X1 port map( A => n3321, ZN => n3147);
   U4547 : INV_X1 port map( A => n3321, ZN => n3148);
   U4548 : INV_X1 port map( A => n3319, ZN => n3150);
   U4549 : INV_X1 port map( A => n3319, ZN => n3151);
   U4550 : INV_X1 port map( A => n3319, ZN => n3152);
   U4551 : INV_X1 port map( A => n3319, ZN => n3154);
   U4552 : INV_X1 port map( A => n3319, ZN => n3155);
   U4553 : INV_X1 port map( A => n3319, ZN => n3156);
   U4554 : INV_X1 port map( A => n3319, ZN => n3158);
   U4555 : INV_X1 port map( A => n3318, ZN => n3159);
   U4556 : INV_X1 port map( A => n3318, ZN => n3160);
   U4557 : INV_X1 port map( A => n3318, ZN => n3162);
   U4558 : INV_X1 port map( A => n3318, ZN => n3163);
   U4559 : INV_X1 port map( A => n3318, ZN => n3164);
   U4560 : INV_X1 port map( A => n3318, ZN => n3166);
   U4561 : INV_X1 port map( A => n3317, ZN => n3167);
   U4562 : INV_X1 port map( A => n3317, ZN => n3168);
   U4563 : INV_X1 port map( A => n3317, ZN => n3170);
   U4564 : INV_X1 port map( A => n3317, ZN => n3171);
   U4565 : INV_X1 port map( A => n3317, ZN => n3172);
   U4566 : INV_X1 port map( A => n3317, ZN => n3174);
   U4567 : INV_X1 port map( A => n3317, ZN => n3175);
   U4568 : INV_X1 port map( A => n3315, ZN => n3176);
   U4569 : INV_X1 port map( A => n3315, ZN => n3178);
   U4570 : INV_X1 port map( A => n3315, ZN => n3180);
   U4571 : INV_X1 port map( A => n3315, ZN => n3181);
   U4572 : INV_X1 port map( A => n3315, ZN => n3183);
   U4573 : INV_X1 port map( A => n3315, ZN => n3184);
   U4574 : INV_X1 port map( A => n3315, ZN => n3185);
   U4575 : INV_X1 port map( A => n3314, ZN => n3187);
   U4576 : INV_X1 port map( A => n3314, ZN => n3188);
   U4577 : INV_X1 port map( A => n3314, ZN => n3189);
   U4578 : INV_X1 port map( A => n3314, ZN => n3191);
   U4579 : INV_X1 port map( A => n3314, ZN => n3192);
   U4580 : INV_X1 port map( A => n3314, ZN => n3193);
   U4581 : INV_X1 port map( A => n3314, ZN => n3195);
   U4582 : INV_X1 port map( A => n3313, ZN => n3196);
   U4583 : INV_X1 port map( A => n3313, ZN => n3197);
   U4584 : INV_X1 port map( A => n3313, ZN => n3199);
   U4585 : INV_X1 port map( A => n3313, ZN => n3200);
   U4586 : INV_X1 port map( A => n3313, ZN => n3201);
   U4587 : INV_X1 port map( A => n3313, ZN => n3203);
   U4588 : INV_X1 port map( A => n3313, ZN => n3204);
   U4589 : INV_X1 port map( A => n3311, ZN => n3205);
   U4590 : INV_X1 port map( A => n3311, ZN => n3207);
   U4591 : INV_X1 port map( A => n3311, ZN => n3208);
   U4592 : INV_X1 port map( A => n3311, ZN => n3209);
   U4593 : INV_X1 port map( A => n3311, ZN => n3211);
   U4594 : INV_X1 port map( A => n3311, ZN => n3212);
   U4595 : INV_X1 port map( A => n3311, ZN => n3213);
   U4596 : INV_X1 port map( A => n3310, ZN => n3215);
   U4597 : INV_X1 port map( A => n3310, ZN => n3216);
   U4598 : INV_X1 port map( A => n3310, ZN => n3217);
   U4599 : INV_X1 port map( A => n3310, ZN => n3219);
   U4600 : INV_X1 port map( A => n3310, ZN => n3220);
   U4601 : INV_X1 port map( A => n3310, ZN => n3221);
   U4602 : INV_X1 port map( A => n3310, ZN => n3223);
   U4603 : INV_X1 port map( A => n3308, ZN => n3224);
   U4604 : INV_X1 port map( A => n3308, ZN => n3225);
   U4605 : INV_X1 port map( A => n3308, ZN => n3227);
   U4606 : INV_X1 port map( A => n3308, ZN => n3228);
   U4607 : INV_X1 port map( A => n3308, ZN => n3229);
   U4608 : INV_X1 port map( A => n3308, ZN => n3231);
   U4609 : INV_X1 port map( A => n3308, ZN => n3232);
   U4610 : INV_X1 port map( A => n3306, ZN => n3233);
   U4611 : INV_X1 port map( A => n3306, ZN => n3235);
   U4612 : INV_X1 port map( A => n3306, ZN => n3236);
   U4613 : INV_X1 port map( A => n3306, ZN => n3237);
   U4614 : INV_X1 port map( A => n3306, ZN => n3239);
   U4615 : INV_X1 port map( A => n3306, ZN => n3240);
   U4616 : INV_X1 port map( A => n3306, ZN => n3241);
   U4617 : INV_X1 port map( A => n3305, ZN => n3243);
   U4618 : INV_X1 port map( A => n3305, ZN => n3245);
   U4619 : INV_X1 port map( A => n3305, ZN => n3246);
   U4620 : INV_X1 port map( A => n3305, ZN => n3248);
   U4621 : INV_X1 port map( A => n3305, ZN => n3249);
   U4622 : INV_X1 port map( A => n3305, ZN => n3250);
   U4623 : INV_X1 port map( A => n3305, ZN => n3252);
   U4624 : INV_X1 port map( A => n3304, ZN => n3253);
   U4625 : INV_X1 port map( A => n3304, ZN => n3254);
   U4626 : INV_X1 port map( A => n3304, ZN => n3256);
   U4627 : INV_X1 port map( A => n3304, ZN => n3257);
   U4628 : INV_X1 port map( A => n3304, ZN => n3258);
   U4629 : INV_X1 port map( A => n3304, ZN => n3260);
   U4630 : INV_X1 port map( A => n3304, ZN => n3261);
   U4631 : INV_X1 port map( A => n3318, ZN => n3262);
   U4632 : INV_X1 port map( A => n3286, ZN => n3264);
   U4633 : NAND2_X1 port map( A1 => ADD_WR(4), A2 => ADD_WR(3), ZN => N2151);
   U4634 : NAND2_X1 port map( A1 => ADD_RD1(4), A2 => ADD_RD1(3), ZN => N8415);
   U4635 : NAND2_X1 port map( A1 => ADD_RD2(4), A2 => ADD_RD2(3), ZN => N8559);
   U4636 : MUX2_X1 port map( A => REGISTERS_87_31_port, B => n2947, S => n1431,
                           Z => n9101);
   U4637 : MUX2_X1 port map( A => REGISTERS_87_30_port, B => n2936, S => n1431,
                           Z => n9102);
   U4638 : MUX2_X1 port map( A => REGISTERS_87_29_port, B => n2925, S => n1431,
                           Z => n9103);
   U4639 : MUX2_X1 port map( A => REGISTERS_87_28_port, B => n2909, S => n1431,
                           Z => n9104);
   U4640 : MUX2_X1 port map( A => REGISTERS_87_27_port, B => n2897, S => n1431,
                           Z => n9105);
   U4641 : MUX2_X1 port map( A => REGISTERS_87_26_port, B => n2886, S => n1431,
                           Z => n9106);
   U4642 : MUX2_X1 port map( A => REGISTERS_87_25_port, B => n2875, S => n1431,
                           Z => n9107);
   U4643 : MUX2_X1 port map( A => REGISTERS_87_24_port, B => n2864, S => n1431,
                           Z => n9108);
   U4644 : MUX2_X1 port map( A => REGISTERS_87_23_port, B => n2853, S => n1431,
                           Z => n9109);
   U4645 : MUX2_X1 port map( A => REGISTERS_87_22_port, B => n2842, S => n1431,
                           Z => n9110);
   U4646 : MUX2_X1 port map( A => REGISTERS_87_21_port, B => n2831, S => n1431,
                           Z => n9111);
   U4647 : MUX2_X1 port map( A => REGISTERS_87_20_port, B => n2820, S => n1431,
                           Z => n9112);
   U4648 : MUX2_X1 port map( A => REGISTERS_87_19_port, B => n2809, S => n1432,
                           Z => n9113);
   U4649 : MUX2_X1 port map( A => REGISTERS_87_18_port, B => n2798, S => n1432,
                           Z => n9114);
   U4650 : MUX2_X1 port map( A => REGISTERS_87_17_port, B => n2787, S => n1432,
                           Z => n9115);
   U4651 : MUX2_X1 port map( A => REGISTERS_87_16_port, B => n2776, S => n1432,
                           Z => n9116);
   U4652 : MUX2_X1 port map( A => REGISTERS_87_15_port, B => n2765, S => n1432,
                           Z => n9117);
   U4653 : MUX2_X1 port map( A => REGISTERS_87_14_port, B => n2754, S => n1432,
                           Z => n9118);
   U4654 : MUX2_X1 port map( A => REGISTERS_87_13_port, B => n2743, S => n1432,
                           Z => n9119);
   U4655 : MUX2_X1 port map( A => REGISTERS_87_12_port, B => n2732, S => n1432,
                           Z => n9120);
   U4656 : MUX2_X1 port map( A => REGISTERS_87_11_port, B => n2721, S => n1432,
                           Z => n9121);
   U4657 : MUX2_X1 port map( A => REGISTERS_87_10_port, B => n2710, S => n1432,
                           Z => n9122);
   U4658 : MUX2_X1 port map( A => REGISTERS_87_9_port, B => n2603, S => n1432, 
                           Z => n9123);
   U4659 : MUX2_X1 port map( A => REGISTERS_87_8_port, B => n2592, S => n1432, 
                           Z => n9124);
   U4660 : MUX2_X1 port map( A => REGISTERS_87_7_port, B => n2581, S => n1433, 
                           Z => n9125);
   U4661 : MUX2_X1 port map( A => REGISTERS_87_6_port, B => n2570, S => n1433, 
                           Z => n9126);
   U4662 : MUX2_X1 port map( A => REGISTERS_87_5_port, B => n2559, S => n1433, 
                           Z => n9127);
   U4663 : MUX2_X1 port map( A => REGISTERS_87_4_port, B => n2548, S => n1433, 
                           Z => n9128);
   U4664 : MUX2_X1 port map( A => REGISTERS_87_3_port, B => n1833, S => n1433, 
                           Z => n9129);
   U4665 : MUX2_X1 port map( A => REGISTERS_87_2_port, B => n1822, S => n1433, 
                           Z => n9130);
   U4666 : MUX2_X1 port map( A => REGISTERS_87_1_port, B => n1811, S => n1433, 
                           Z => n9131);
   U4667 : MUX2_X1 port map( A => REGISTERS_87_0_port, B => n1800, S => n1433, 
                           Z => n9132);
   U4668 : MUX2_X1 port map( A => REGISTERS_86_31_port, B => n2947, S => n1434,
                           Z => n9069);
   U4669 : MUX2_X1 port map( A => REGISTERS_86_30_port, B => n2936, S => n1434,
                           Z => n9070);
   U4670 : MUX2_X1 port map( A => REGISTERS_86_29_port, B => n2925, S => n1434,
                           Z => n9071);
   U4671 : MUX2_X1 port map( A => REGISTERS_86_28_port, B => n2909, S => n1434,
                           Z => n9072);
   U4672 : MUX2_X1 port map( A => REGISTERS_86_27_port, B => n2897, S => n1434,
                           Z => n9073);
   U4673 : MUX2_X1 port map( A => REGISTERS_86_26_port, B => n2886, S => n1434,
                           Z => n9074);
   U4674 : MUX2_X1 port map( A => REGISTERS_86_25_port, B => n2875, S => n1434,
                           Z => n9075);
   U4675 : MUX2_X1 port map( A => REGISTERS_86_24_port, B => n2864, S => n1434,
                           Z => n9076);
   U4676 : MUX2_X1 port map( A => REGISTERS_86_23_port, B => n2853, S => n1434,
                           Z => n9077);
   U4677 : MUX2_X1 port map( A => REGISTERS_86_22_port, B => n2842, S => n1434,
                           Z => n9078);
   U4678 : MUX2_X1 port map( A => REGISTERS_86_21_port, B => n2831, S => n1434,
                           Z => n9079);
   U4679 : MUX2_X1 port map( A => REGISTERS_86_20_port, B => n2820, S => n1434,
                           Z => n9080);
   U4680 : MUX2_X1 port map( A => REGISTERS_86_19_port, B => n2809, S => n1435,
                           Z => n9081);
   U4681 : MUX2_X1 port map( A => REGISTERS_86_18_port, B => n2798, S => n1435,
                           Z => n9082);
   U4682 : MUX2_X1 port map( A => REGISTERS_86_17_port, B => n2787, S => n1435,
                           Z => n9083);
   U4683 : MUX2_X1 port map( A => REGISTERS_86_16_port, B => n2776, S => n1435,
                           Z => n9084);
   U4684 : MUX2_X1 port map( A => REGISTERS_86_15_port, B => n2765, S => n1435,
                           Z => n9085);
   U4685 : MUX2_X1 port map( A => REGISTERS_86_14_port, B => n2754, S => n1435,
                           Z => n9086);
   U4686 : MUX2_X1 port map( A => REGISTERS_86_13_port, B => n2743, S => n1435,
                           Z => n9087);
   U4687 : MUX2_X1 port map( A => REGISTERS_86_12_port, B => n2732, S => n1435,
                           Z => n9088);
   U4688 : MUX2_X1 port map( A => REGISTERS_86_11_port, B => n2721, S => n1435,
                           Z => n9089);
   U4689 : MUX2_X1 port map( A => REGISTERS_86_10_port, B => n2710, S => n1435,
                           Z => n9090);
   U4690 : MUX2_X1 port map( A => REGISTERS_86_9_port, B => n2603, S => n1435, 
                           Z => n9091);
   U4691 : MUX2_X1 port map( A => REGISTERS_86_8_port, B => n2592, S => n1435, 
                           Z => n9092);
   U4692 : MUX2_X1 port map( A => REGISTERS_86_7_port, B => n2581, S => n1436, 
                           Z => n9093);
   U4693 : MUX2_X1 port map( A => REGISTERS_86_6_port, B => n2570, S => n1436, 
                           Z => n9094);
   U4694 : MUX2_X1 port map( A => REGISTERS_86_5_port, B => n2559, S => n1436, 
                           Z => n9095);
   U4695 : MUX2_X1 port map( A => REGISTERS_86_4_port, B => n2548, S => n1436, 
                           Z => n9096);
   U4696 : MUX2_X1 port map( A => REGISTERS_86_3_port, B => n1833, S => n1436, 
                           Z => n9097);
   U4697 : MUX2_X1 port map( A => REGISTERS_86_2_port, B => n1822, S => n1436, 
                           Z => n9098);
   U4698 : MUX2_X1 port map( A => REGISTERS_86_1_port, B => n1811, S => n1436, 
                           Z => n9099);
   U4699 : MUX2_X1 port map( A => REGISTERS_86_0_port, B => n1800, S => n1436, 
                           Z => n9100);
   U4700 : MUX2_X1 port map( A => REGISTERS_85_31_port, B => n2947, S => n1437,
                           Z => n9037);
   U4701 : MUX2_X1 port map( A => REGISTERS_85_30_port, B => n2936, S => n1437,
                           Z => n9038);
   U4702 : MUX2_X1 port map( A => REGISTERS_85_29_port, B => n2925, S => n1437,
                           Z => n9039);
   U4703 : MUX2_X1 port map( A => REGISTERS_85_28_port, B => n2909, S => n1437,
                           Z => n9040);
   U4704 : MUX2_X1 port map( A => REGISTERS_85_27_port, B => n2897, S => n1437,
                           Z => n9041);
   U4705 : MUX2_X1 port map( A => REGISTERS_85_26_port, B => n2886, S => n1437,
                           Z => n9042);
   U4706 : MUX2_X1 port map( A => REGISTERS_85_25_port, B => n2875, S => n1437,
                           Z => n9043);
   U4707 : MUX2_X1 port map( A => REGISTERS_85_24_port, B => n2864, S => n1437,
                           Z => n9044);
   U4708 : MUX2_X1 port map( A => REGISTERS_85_23_port, B => n2853, S => n1437,
                           Z => n9045);
   U4709 : MUX2_X1 port map( A => REGISTERS_85_22_port, B => n2842, S => n1437,
                           Z => n9046);
   U4710 : MUX2_X1 port map( A => REGISTERS_85_21_port, B => n2831, S => n1437,
                           Z => n9047);
   U4711 : MUX2_X1 port map( A => REGISTERS_85_20_port, B => n2820, S => n1437,
                           Z => n9048);
   U4712 : MUX2_X1 port map( A => REGISTERS_85_19_port, B => n2809, S => n1438,
                           Z => n9049);
   U4713 : MUX2_X1 port map( A => REGISTERS_85_18_port, B => n2798, S => n1438,
                           Z => n9050);
   U4714 : MUX2_X1 port map( A => REGISTERS_85_17_port, B => n2787, S => n1438,
                           Z => n9051);
   U4715 : MUX2_X1 port map( A => REGISTERS_85_16_port, B => n2776, S => n1438,
                           Z => n9052);
   U4716 : MUX2_X1 port map( A => REGISTERS_85_15_port, B => n2765, S => n1438,
                           Z => n9053);
   U4717 : MUX2_X1 port map( A => REGISTERS_85_14_port, B => n2754, S => n1438,
                           Z => n9054);
   U4718 : MUX2_X1 port map( A => REGISTERS_85_13_port, B => n2743, S => n1438,
                           Z => n9055);
   U4719 : MUX2_X1 port map( A => REGISTERS_85_12_port, B => n2732, S => n1438,
                           Z => n9056);
   U4720 : MUX2_X1 port map( A => REGISTERS_85_11_port, B => n2721, S => n1438,
                           Z => n9057);
   U4721 : MUX2_X1 port map( A => REGISTERS_85_10_port, B => n2710, S => n1438,
                           Z => n9058);
   U4722 : MUX2_X1 port map( A => REGISTERS_85_9_port, B => n2603, S => n1438, 
                           Z => n9059);
   U4723 : MUX2_X1 port map( A => REGISTERS_85_8_port, B => n2592, S => n1438, 
                           Z => n9060);
   U4724 : MUX2_X1 port map( A => REGISTERS_85_7_port, B => n2581, S => n1439, 
                           Z => n9061);
   U4725 : MUX2_X1 port map( A => REGISTERS_85_6_port, B => n2570, S => n1439, 
                           Z => n9062);
   U4726 : MUX2_X1 port map( A => REGISTERS_85_5_port, B => n2559, S => n1439, 
                           Z => n9063);
   U4727 : MUX2_X1 port map( A => REGISTERS_85_4_port, B => n2548, S => n1439, 
                           Z => n9064);
   U4728 : MUX2_X1 port map( A => REGISTERS_85_3_port, B => n1833, S => n1439, 
                           Z => n9065);
   U4729 : MUX2_X1 port map( A => REGISTERS_85_2_port, B => n1822, S => n1439, 
                           Z => n9066);
   U4730 : MUX2_X1 port map( A => REGISTERS_85_1_port, B => n1811, S => n1439, 
                           Z => n9067);
   U4731 : MUX2_X1 port map( A => REGISTERS_85_0_port, B => n1800, S => n1439, 
                           Z => n9068);
   U4732 : MUX2_X1 port map( A => REGISTERS_84_31_port, B => n2947, S => n1440,
                           Z => n9005);
   U4733 : MUX2_X1 port map( A => REGISTERS_84_30_port, B => n2936, S => n1440,
                           Z => n9006);
   U4734 : MUX2_X1 port map( A => REGISTERS_84_29_port, B => n2925, S => n1440,
                           Z => n9007);
   U4735 : MUX2_X1 port map( A => REGISTERS_84_28_port, B => n2909, S => n1440,
                           Z => n9008);
   U4736 : MUX2_X1 port map( A => REGISTERS_84_27_port, B => n2897, S => n1440,
                           Z => n9009);
   U4737 : MUX2_X1 port map( A => REGISTERS_84_26_port, B => n2886, S => n1440,
                           Z => n9010);
   U4738 : MUX2_X1 port map( A => REGISTERS_84_25_port, B => n2875, S => n1440,
                           Z => n9011);
   U4739 : MUX2_X1 port map( A => REGISTERS_84_24_port, B => n2864, S => n1440,
                           Z => n9012);
   U4740 : MUX2_X1 port map( A => REGISTERS_84_23_port, B => n2853, S => n1440,
                           Z => n9013);
   U4741 : MUX2_X1 port map( A => REGISTERS_84_22_port, B => n2842, S => n1440,
                           Z => n9014);
   U4742 : MUX2_X1 port map( A => REGISTERS_84_21_port, B => n2831, S => n1440,
                           Z => n9015);
   U4743 : MUX2_X1 port map( A => REGISTERS_84_20_port, B => n2820, S => n1440,
                           Z => n9016);
   U4744 : MUX2_X1 port map( A => REGISTERS_84_19_port, B => n2809, S => n1441,
                           Z => n9017);
   U4745 : MUX2_X1 port map( A => REGISTERS_84_18_port, B => n2798, S => n1441,
                           Z => n9018);
   U4746 : MUX2_X1 port map( A => REGISTERS_84_17_port, B => n2787, S => n1441,
                           Z => n9019);
   U4747 : MUX2_X1 port map( A => REGISTERS_84_16_port, B => n2776, S => n1441,
                           Z => n9020);
   U4748 : MUX2_X1 port map( A => REGISTERS_84_15_port, B => n2765, S => n1441,
                           Z => n9021);
   U4749 : MUX2_X1 port map( A => REGISTERS_84_14_port, B => n2754, S => n1441,
                           Z => n9022);
   U4750 : MUX2_X1 port map( A => REGISTERS_84_13_port, B => n2743, S => n1441,
                           Z => n9023);
   U4751 : MUX2_X1 port map( A => REGISTERS_84_12_port, B => n2732, S => n1441,
                           Z => n9024);
   U4752 : MUX2_X1 port map( A => REGISTERS_84_11_port, B => n2721, S => n1441,
                           Z => n9025);
   U4753 : MUX2_X1 port map( A => REGISTERS_84_10_port, B => n2710, S => n1441,
                           Z => n9026);
   U4754 : MUX2_X1 port map( A => REGISTERS_84_9_port, B => n2603, S => n1441, 
                           Z => n9027);
   U4755 : MUX2_X1 port map( A => REGISTERS_84_8_port, B => n2592, S => n1441, 
                           Z => n9028);
   U4756 : MUX2_X1 port map( A => REGISTERS_84_7_port, B => n2581, S => n1442, 
                           Z => n9029);
   U4757 : MUX2_X1 port map( A => REGISTERS_84_6_port, B => n2570, S => n1442, 
                           Z => n9030);
   U4758 : MUX2_X1 port map( A => REGISTERS_84_5_port, B => n2559, S => n1442, 
                           Z => n9031);
   U4759 : MUX2_X1 port map( A => REGISTERS_84_4_port, B => n2548, S => n1442, 
                           Z => n9032);
   U4760 : MUX2_X1 port map( A => REGISTERS_84_3_port, B => n1833, S => n1442, 
                           Z => n9033);
   U4761 : MUX2_X1 port map( A => REGISTERS_84_2_port, B => n1822, S => n1442, 
                           Z => n9034);
   U4762 : MUX2_X1 port map( A => REGISTERS_84_1_port, B => n1811, S => n1442, 
                           Z => n9035);
   U4763 : MUX2_X1 port map( A => REGISTERS_84_0_port, B => n1800, S => n1442, 
                           Z => n9036);
   U4764 : MUX2_X1 port map( A => REGISTERS_83_31_port, B => n2947, S => n1443,
                           Z => n8973);
   U4765 : MUX2_X1 port map( A => REGISTERS_83_30_port, B => n2936, S => n1443,
                           Z => n8974);
   U4766 : MUX2_X1 port map( A => REGISTERS_83_29_port, B => n2925, S => n1443,
                           Z => n8975);
   U4767 : MUX2_X1 port map( A => REGISTERS_83_28_port, B => n2909, S => n1443,
                           Z => n8976);
   U4768 : MUX2_X1 port map( A => REGISTERS_83_27_port, B => n2897, S => n1443,
                           Z => n8977);
   U4769 : MUX2_X1 port map( A => REGISTERS_83_26_port, B => n2886, S => n1443,
                           Z => n8978);
   U4770 : MUX2_X1 port map( A => REGISTERS_83_25_port, B => n2875, S => n1443,
                           Z => n8979);
   U4771 : MUX2_X1 port map( A => REGISTERS_83_24_port, B => n2864, S => n1443,
                           Z => n8980);
   U4772 : MUX2_X1 port map( A => REGISTERS_83_23_port, B => n2853, S => n1443,
                           Z => n8981);
   U4773 : MUX2_X1 port map( A => REGISTERS_83_22_port, B => n2842, S => n1443,
                           Z => n8982);
   U4774 : MUX2_X1 port map( A => REGISTERS_83_21_port, B => n2831, S => n1443,
                           Z => n8983);
   U4775 : MUX2_X1 port map( A => REGISTERS_83_20_port, B => n2820, S => n1443,
                           Z => n8984);
   U4776 : MUX2_X1 port map( A => REGISTERS_83_19_port, B => n2809, S => n1444,
                           Z => n8985);
   U4777 : MUX2_X1 port map( A => REGISTERS_83_18_port, B => n2798, S => n1444,
                           Z => n8986);
   U4778 : MUX2_X1 port map( A => REGISTERS_83_17_port, B => n2787, S => n1444,
                           Z => n8987);
   U4779 : MUX2_X1 port map( A => REGISTERS_83_16_port, B => n2776, S => n1444,
                           Z => n8988);
   U4780 : MUX2_X1 port map( A => REGISTERS_83_15_port, B => n2765, S => n1444,
                           Z => n8989);
   U4781 : MUX2_X1 port map( A => REGISTERS_83_14_port, B => n2754, S => n1444,
                           Z => n8990);
   U4782 : MUX2_X1 port map( A => REGISTERS_83_13_port, B => n2743, S => n1444,
                           Z => n8991);
   U4783 : MUX2_X1 port map( A => REGISTERS_83_12_port, B => n2732, S => n1444,
                           Z => n8992);
   U4784 : MUX2_X1 port map( A => REGISTERS_83_11_port, B => n2721, S => n1444,
                           Z => n8993);
   U4785 : MUX2_X1 port map( A => REGISTERS_83_10_port, B => n2710, S => n1444,
                           Z => n8994);
   U4786 : MUX2_X1 port map( A => REGISTERS_83_9_port, B => n2603, S => n1444, 
                           Z => n8995);
   U4787 : MUX2_X1 port map( A => REGISTERS_83_8_port, B => n2592, S => n1444, 
                           Z => n8996);
   U4788 : MUX2_X1 port map( A => REGISTERS_83_7_port, B => n2581, S => n1445, 
                           Z => n8997);
   U4789 : MUX2_X1 port map( A => REGISTERS_83_6_port, B => n2570, S => n1445, 
                           Z => n8998);
   U4790 : MUX2_X1 port map( A => REGISTERS_83_5_port, B => n2559, S => n1445, 
                           Z => n8999);
   U4791 : MUX2_X1 port map( A => REGISTERS_83_4_port, B => n2548, S => n1445, 
                           Z => n9000);
   U4792 : MUX2_X1 port map( A => REGISTERS_83_3_port, B => n1833, S => n1445, 
                           Z => n9001);
   U4793 : MUX2_X1 port map( A => REGISTERS_83_2_port, B => n1822, S => n1445, 
                           Z => n9002);
   U4794 : MUX2_X1 port map( A => REGISTERS_83_1_port, B => n1811, S => n1445, 
                           Z => n9003);
   U4795 : MUX2_X1 port map( A => REGISTERS_83_0_port, B => n1800, S => n1445, 
                           Z => n9004);
   U4796 : MUX2_X1 port map( A => REGISTERS_82_31_port, B => n2947, S => n1446,
                           Z => n8941);
   U4797 : MUX2_X1 port map( A => REGISTERS_82_30_port, B => n2936, S => n1446,
                           Z => n8942);
   U4798 : MUX2_X1 port map( A => REGISTERS_82_29_port, B => n2925, S => n1446,
                           Z => n8943);
   U4799 : MUX2_X1 port map( A => REGISTERS_82_28_port, B => n2909, S => n1446,
                           Z => n8944);
   U4800 : MUX2_X1 port map( A => REGISTERS_82_27_port, B => n2897, S => n1446,
                           Z => n8945);
   U4801 : MUX2_X1 port map( A => REGISTERS_82_26_port, B => n2886, S => n1446,
                           Z => n8946);
   U4802 : MUX2_X1 port map( A => REGISTERS_82_25_port, B => n2875, S => n1446,
                           Z => n8947);
   U4803 : MUX2_X1 port map( A => REGISTERS_82_24_port, B => n2864, S => n1446,
                           Z => n8948);
   U4804 : MUX2_X1 port map( A => REGISTERS_82_23_port, B => n2853, S => n1446,
                           Z => n8949);
   U4805 : MUX2_X1 port map( A => REGISTERS_82_22_port, B => n2842, S => n1446,
                           Z => n8950);
   U4806 : MUX2_X1 port map( A => REGISTERS_82_21_port, B => n2831, S => n1446,
                           Z => n8951);
   U4807 : MUX2_X1 port map( A => REGISTERS_82_20_port, B => n2820, S => n1446,
                           Z => n8952);
   U4808 : MUX2_X1 port map( A => REGISTERS_82_19_port, B => n2809, S => n1447,
                           Z => n8953);
   U4809 : MUX2_X1 port map( A => REGISTERS_82_18_port, B => n2798, S => n1447,
                           Z => n8954);
   U4810 : MUX2_X1 port map( A => REGISTERS_82_17_port, B => n2787, S => n1447,
                           Z => n8955);
   U4811 : MUX2_X1 port map( A => REGISTERS_82_16_port, B => n2776, S => n1447,
                           Z => n8956);
   U4812 : MUX2_X1 port map( A => REGISTERS_82_15_port, B => n2765, S => n1447,
                           Z => n8957);
   U4813 : MUX2_X1 port map( A => REGISTERS_82_14_port, B => n2754, S => n1447,
                           Z => n8958);
   U4814 : MUX2_X1 port map( A => REGISTERS_82_13_port, B => n2743, S => n1447,
                           Z => n8959);
   U4815 : MUX2_X1 port map( A => REGISTERS_82_12_port, B => n2732, S => n1447,
                           Z => n8960);
   U4816 : MUX2_X1 port map( A => REGISTERS_82_11_port, B => n2721, S => n1447,
                           Z => n8961);
   U4817 : MUX2_X1 port map( A => REGISTERS_82_10_port, B => n2710, S => n1447,
                           Z => n8962);
   U4818 : MUX2_X1 port map( A => REGISTERS_82_9_port, B => n2603, S => n1447, 
                           Z => n8963);
   U4819 : MUX2_X1 port map( A => REGISTERS_82_8_port, B => n2592, S => n1447, 
                           Z => n8964);
   U4820 : MUX2_X1 port map( A => REGISTERS_82_7_port, B => n2581, S => n1448, 
                           Z => n8965);
   U4821 : MUX2_X1 port map( A => REGISTERS_82_6_port, B => n2570, S => n1448, 
                           Z => n8966);
   U4822 : MUX2_X1 port map( A => REGISTERS_82_5_port, B => n2559, S => n1448, 
                           Z => n8967);
   U4823 : MUX2_X1 port map( A => REGISTERS_82_4_port, B => n2548, S => n1448, 
                           Z => n8968);
   U4824 : MUX2_X1 port map( A => REGISTERS_82_3_port, B => n1833, S => n1448, 
                           Z => n8969);
   U4825 : MUX2_X1 port map( A => REGISTERS_82_2_port, B => n1822, S => n1448, 
                           Z => n8970);
   U4826 : MUX2_X1 port map( A => REGISTERS_82_1_port, B => n1811, S => n1448, 
                           Z => n8971);
   U4827 : MUX2_X1 port map( A => REGISTERS_82_0_port, B => n1800, S => n1448, 
                           Z => n8972);
   U4828 : MUX2_X1 port map( A => n10886, B => n2947, S => n1449, Z => n8909);
   U4829 : MUX2_X1 port map( A => n10887, B => n2936, S => n1449, Z => n8910);
   U4830 : MUX2_X1 port map( A => n10888, B => n2925, S => n1449, Z => n8911);
   U4831 : MUX2_X1 port map( A => n10889, B => n2909, S => n1449, Z => n8912);
   U4832 : MUX2_X1 port map( A => n10890, B => n2897, S => n1449, Z => n8913);
   U4833 : MUX2_X1 port map( A => n10891, B => n2886, S => n1449, Z => n8914);
   U4834 : MUX2_X1 port map( A => n10892, B => n2875, S => n1449, Z => n8915);
   U4835 : MUX2_X1 port map( A => n10893, B => n2864, S => n1449, Z => n8916);
   U4836 : MUX2_X1 port map( A => n10894, B => n2853, S => n1449, Z => n8917);
   U4837 : MUX2_X1 port map( A => n10895, B => n2842, S => n1449, Z => n8918);
   U4838 : MUX2_X1 port map( A => n10896, B => n2831, S => n1449, Z => n8919);
   U4839 : MUX2_X1 port map( A => n10897, B => n2820, S => n1449, Z => n8920);
   U4840 : MUX2_X1 port map( A => n10898, B => n2809, S => n1450, Z => n8921);
   U4841 : MUX2_X1 port map( A => n10899, B => n2798, S => n1450, Z => n8922);
   U4842 : MUX2_X1 port map( A => n10900, B => n2787, S => n1450, Z => n8923);
   U4843 : MUX2_X1 port map( A => n10901, B => n2776, S => n1450, Z => n8924);
   U4844 : MUX2_X1 port map( A => n10902, B => n2765, S => n1450, Z => n8925);
   U4845 : MUX2_X1 port map( A => n10903, B => n2754, S => n1450, Z => n8926);
   U4846 : MUX2_X1 port map( A => n10904, B => n2743, S => n1450, Z => n8927);
   U4847 : MUX2_X1 port map( A => n10905, B => n2732, S => n1450, Z => n8928);
   U4848 : MUX2_X1 port map( A => n10906, B => n2721, S => n1450, Z => n8929);
   U4849 : MUX2_X1 port map( A => n10907, B => n2710, S => n1450, Z => n8930);
   U4850 : MUX2_X1 port map( A => n10908, B => n2603, S => n1450, Z => n8931);
   U4851 : MUX2_X1 port map( A => n10909, B => n2592, S => n1450, Z => n8932);
   U4852 : MUX2_X1 port map( A => n10910, B => n2581, S => n1451, Z => n8933);
   U4853 : MUX2_X1 port map( A => n10911, B => n2570, S => n1451, Z => n8934);
   U4854 : MUX2_X1 port map( A => n10912, B => n2559, S => n1451, Z => n8935);
   U4855 : MUX2_X1 port map( A => n10913, B => n2548, S => n1451, Z => n8936);
   U4856 : MUX2_X1 port map( A => n10914, B => n1833, S => n1451, Z => n8937);
   U4857 : MUX2_X1 port map( A => n10915, B => n1822, S => n1451, Z => n8938);
   U4858 : MUX2_X1 port map( A => n10916, B => n1811, S => n1451, Z => n8939);
   U4859 : MUX2_X1 port map( A => n10917, B => n1800, S => n1451, Z => n8940);
   U4860 : MUX2_X1 port map( A => n10854, B => n2947, S => n1452, Z => n8877);
   U4861 : MUX2_X1 port map( A => n10855, B => n2936, S => n1452, Z => n8878);
   U4862 : MUX2_X1 port map( A => n10856, B => n2925, S => n1452, Z => n8879);
   U4863 : MUX2_X1 port map( A => n10857, B => n2909, S => n1452, Z => n8880);
   U4864 : MUX2_X1 port map( A => n10858, B => n2897, S => n1452, Z => n8881);
   U4865 : MUX2_X1 port map( A => n10859, B => n2886, S => n1452, Z => n8882);
   U4866 : MUX2_X1 port map( A => n10860, B => n2875, S => n1452, Z => n8883);
   U4867 : MUX2_X1 port map( A => n10861, B => n2864, S => n1452, Z => n8884);
   U4868 : MUX2_X1 port map( A => n10862, B => n2853, S => n1452, Z => n8885);
   U4869 : MUX2_X1 port map( A => n10863, B => n2842, S => n1452, Z => n8886);
   U4870 : MUX2_X1 port map( A => n10864, B => n2831, S => n1452, Z => n8887);
   U4871 : MUX2_X1 port map( A => n10865, B => n2820, S => n1452, Z => n8888);
   U4872 : MUX2_X1 port map( A => n10866, B => n2809, S => n1453, Z => n8889);
   U4873 : MUX2_X1 port map( A => n10867, B => n2798, S => n1453, Z => n8890);
   U4874 : MUX2_X1 port map( A => n10868, B => n2787, S => n1453, Z => n8891);
   U4875 : MUX2_X1 port map( A => n10869, B => n2776, S => n1453, Z => n8892);
   U4876 : MUX2_X1 port map( A => n10870, B => n2765, S => n1453, Z => n8893);
   U4877 : MUX2_X1 port map( A => n10871, B => n2754, S => n1453, Z => n8894);
   U4878 : MUX2_X1 port map( A => n10872, B => n2743, S => n1453, Z => n8895);
   U4879 : MUX2_X1 port map( A => n10873, B => n2732, S => n1453, Z => n8896);
   U4880 : MUX2_X1 port map( A => n10874, B => n2721, S => n1453, Z => n8897);
   U4881 : MUX2_X1 port map( A => n10875, B => n2710, S => n1453, Z => n8898);
   U4882 : MUX2_X1 port map( A => n10876, B => n2603, S => n1453, Z => n8899);
   U4883 : MUX2_X1 port map( A => n10877, B => n2592, S => n1453, Z => n8900);
   U4884 : MUX2_X1 port map( A => n10878, B => n2581, S => n1454, Z => n8901);
   U4885 : MUX2_X1 port map( A => n10879, B => n2570, S => n1454, Z => n8902);
   U4886 : MUX2_X1 port map( A => n10880, B => n2559, S => n1454, Z => n8903);
   U4887 : MUX2_X1 port map( A => n10881, B => n2548, S => n1454, Z => n8904);
   U4888 : MUX2_X1 port map( A => n10882, B => n1833, S => n1454, Z => n8905);
   U4889 : MUX2_X1 port map( A => n10883, B => n1822, S => n1454, Z => n8906);
   U4890 : MUX2_X1 port map( A => n10884, B => n1811, S => n1454, Z => n8907);
   U4891 : MUX2_X1 port map( A => n10885, B => n1800, S => n1454, Z => n8908);
   U4892 : MUX2_X1 port map( A => n10822, B => n2947, S => n1455, Z => n8845);
   U4893 : MUX2_X1 port map( A => n10823, B => n2936, S => n1455, Z => n8846);
   U4894 : MUX2_X1 port map( A => n10824, B => n2925, S => n1455, Z => n8847);
   U4895 : MUX2_X1 port map( A => n10825, B => n2909, S => n1455, Z => n8848);
   U4896 : MUX2_X1 port map( A => n10826, B => n2897, S => n1455, Z => n8849);
   U4897 : MUX2_X1 port map( A => n10827, B => n2886, S => n1455, Z => n8850);
   U4898 : MUX2_X1 port map( A => n10828, B => n2875, S => n1455, Z => n8851);
   U4899 : MUX2_X1 port map( A => n10829, B => n2864, S => n1455, Z => n8852);
   U4900 : MUX2_X1 port map( A => n10830, B => n2853, S => n1455, Z => n8853);
   U4901 : MUX2_X1 port map( A => n10831, B => n2842, S => n1455, Z => n8854);
   U4902 : MUX2_X1 port map( A => n10832, B => n2831, S => n1455, Z => n8855);
   U4903 : MUX2_X1 port map( A => n10833, B => n2820, S => n1455, Z => n8856);
   U4904 : MUX2_X1 port map( A => n10834, B => n2809, S => n1456, Z => n8857);
   U4905 : MUX2_X1 port map( A => n10835, B => n2798, S => n1456, Z => n8858);
   U4906 : MUX2_X1 port map( A => n10836, B => n2787, S => n1456, Z => n8859);
   U4907 : MUX2_X1 port map( A => n10837, B => n2776, S => n1456, Z => n8860);
   U4908 : MUX2_X1 port map( A => n10838, B => n2765, S => n1456, Z => n8861);
   U4909 : MUX2_X1 port map( A => n10839, B => n2754, S => n1456, Z => n8862);
   U4910 : MUX2_X1 port map( A => n10840, B => n2743, S => n1456, Z => n8863);
   U4911 : MUX2_X1 port map( A => n10841, B => n2732, S => n1456, Z => n8864);
   U4912 : MUX2_X1 port map( A => n10842, B => n2721, S => n1456, Z => n8865);
   U4913 : MUX2_X1 port map( A => n10843, B => n2710, S => n1456, Z => n8866);
   U4914 : MUX2_X1 port map( A => n10844, B => n2603, S => n1456, Z => n8867);
   U4915 : MUX2_X1 port map( A => n10845, B => n2592, S => n1456, Z => n8868);
   U4916 : MUX2_X1 port map( A => n10846, B => n2581, S => n1457, Z => n8869);
   U4917 : MUX2_X1 port map( A => n10847, B => n2570, S => n1457, Z => n8870);
   U4918 : MUX2_X1 port map( A => n10848, B => n2559, S => n1457, Z => n8871);
   U4919 : MUX2_X1 port map( A => n10849, B => n2548, S => n1457, Z => n8872);
   U4920 : MUX2_X1 port map( A => n10850, B => n1833, S => n1457, Z => n8873);
   U4921 : MUX2_X1 port map( A => n10851, B => n1822, S => n1457, Z => n8874);
   U4922 : MUX2_X1 port map( A => n10852, B => n1811, S => n1457, Z => n8875);
   U4923 : MUX2_X1 port map( A => n10853, B => n1800, S => n1457, Z => n8876);
   U4924 : MUX2_X1 port map( A => REGISTERS_78_31_port, B => n2947, S => n1458,
                           Z => n8813);
   U4925 : MUX2_X1 port map( A => REGISTERS_78_30_port, B => n2936, S => n1458,
                           Z => n8814);
   U4926 : MUX2_X1 port map( A => REGISTERS_78_29_port, B => n2925, S => n1458,
                           Z => n8815);
   U4927 : MUX2_X1 port map( A => REGISTERS_78_28_port, B => n2909, S => n1458,
                           Z => n8816);
   U4928 : MUX2_X1 port map( A => REGISTERS_78_27_port, B => n2897, S => n1458,
                           Z => n8817);
   U4929 : MUX2_X1 port map( A => REGISTERS_78_26_port, B => n2886, S => n1458,
                           Z => n8818);
   U4930 : MUX2_X1 port map( A => REGISTERS_78_25_port, B => n2875, S => n1458,
                           Z => n8819);
   U4931 : MUX2_X1 port map( A => REGISTERS_78_24_port, B => n2864, S => n1458,
                           Z => n8820);
   U4932 : MUX2_X1 port map( A => REGISTERS_78_23_port, B => n2853, S => n1458,
                           Z => n8821);
   U4933 : MUX2_X1 port map( A => REGISTERS_78_22_port, B => n2842, S => n1458,
                           Z => n8822);
   U4934 : MUX2_X1 port map( A => REGISTERS_78_21_port, B => n2831, S => n1458,
                           Z => n8823);
   U4935 : MUX2_X1 port map( A => REGISTERS_78_20_port, B => n2820, S => n1458,
                           Z => n8824);
   U4936 : MUX2_X1 port map( A => REGISTERS_78_19_port, B => n2809, S => n1459,
                           Z => n8825);
   U4937 : MUX2_X1 port map( A => REGISTERS_78_18_port, B => n2798, S => n1459,
                           Z => n8826);
   U4938 : MUX2_X1 port map( A => REGISTERS_78_17_port, B => n2787, S => n1459,
                           Z => n8827);
   U4939 : MUX2_X1 port map( A => REGISTERS_78_16_port, B => n2776, S => n1459,
                           Z => n8828);
   U4940 : MUX2_X1 port map( A => REGISTERS_78_15_port, B => n2765, S => n1459,
                           Z => n8829);
   U4941 : MUX2_X1 port map( A => REGISTERS_78_14_port, B => n2754, S => n1459,
                           Z => n8830);
   U4942 : MUX2_X1 port map( A => REGISTERS_78_13_port, B => n2743, S => n1459,
                           Z => n8831);
   U4943 : MUX2_X1 port map( A => REGISTERS_78_12_port, B => n2732, S => n1459,
                           Z => n8832);
   U4944 : MUX2_X1 port map( A => REGISTERS_78_11_port, B => n2721, S => n1459,
                           Z => n8833_port);
   U4945 : MUX2_X1 port map( A => REGISTERS_78_10_port, B => n2710, S => n1459,
                           Z => n8834_port);
   U4946 : MUX2_X1 port map( A => REGISTERS_78_9_port, B => n2603, S => n1459, 
                           Z => n8835);
   U4947 : MUX2_X1 port map( A => REGISTERS_78_8_port, B => n2592, S => n1459, 
                           Z => n8836);
   U4948 : MUX2_X1 port map( A => REGISTERS_78_7_port, B => n2581, S => n1460, 
                           Z => n8837);
   U4949 : MUX2_X1 port map( A => REGISTERS_78_6_port, B => n2570, S => n1460, 
                           Z => n8838);
   U4950 : MUX2_X1 port map( A => REGISTERS_78_5_port, B => n2559, S => n1460, 
                           Z => n8839);
   U4951 : MUX2_X1 port map( A => REGISTERS_78_4_port, B => n2548, S => n1460, 
                           Z => n8840);
   U4952 : MUX2_X1 port map( A => REGISTERS_78_3_port, B => n1833, S => n1460, 
                           Z => n8841);
   U4953 : MUX2_X1 port map( A => REGISTERS_78_2_port, B => n1822, S => n1460, 
                           Z => n8842);
   U4954 : MUX2_X1 port map( A => REGISTERS_78_1_port, B => n1811, S => n1460, 
                           Z => n8843);
   U4955 : MUX2_X1 port map( A => REGISTERS_78_0_port, B => n1800, S => n1460, 
                           Z => n8844);
   U4956 : MUX2_X1 port map( A => REGISTERS_77_31_port, B => n2947, S => n1461,
                           Z => n8781);
   U4957 : MUX2_X1 port map( A => REGISTERS_77_30_port, B => n2936, S => n1461,
                           Z => n8782);
   U4958 : MUX2_X1 port map( A => REGISTERS_77_29_port, B => n2925, S => n1461,
                           Z => n8783);
   U4959 : MUX2_X1 port map( A => REGISTERS_77_28_port, B => n2909, S => n1461,
                           Z => n8784);
   U4960 : MUX2_X1 port map( A => REGISTERS_77_27_port, B => n2897, S => n1461,
                           Z => n8785);
   U4961 : MUX2_X1 port map( A => REGISTERS_77_26_port, B => n2886, S => n1461,
                           Z => n8786);
   U4962 : MUX2_X1 port map( A => REGISTERS_77_25_port, B => n2875, S => n1461,
                           Z => n8787_port);
   U4963 : MUX2_X1 port map( A => REGISTERS_77_24_port, B => n2864, S => n1461,
                           Z => n8788_port);
   U4964 : MUX2_X1 port map( A => REGISTERS_77_23_port, B => n2853, S => n1461,
                           Z => n8789_port);
   U4965 : MUX2_X1 port map( A => REGISTERS_77_22_port, B => n2842, S => n1461,
                           Z => n8790_port);
   U4966 : MUX2_X1 port map( A => REGISTERS_77_21_port, B => n2831, S => n1461,
                           Z => n8791_port);
   U4967 : MUX2_X1 port map( A => REGISTERS_77_20_port, B => n2820, S => n1461,
                           Z => n8792);
   U4968 : MUX2_X1 port map( A => REGISTERS_77_19_port, B => n2809, S => n1462,
                           Z => n8793);
   U4969 : MUX2_X1 port map( A => REGISTERS_77_18_port, B => n2798, S => n1462,
                           Z => n8794);
   U4970 : MUX2_X1 port map( A => REGISTERS_77_17_port, B => n2787, S => n1462,
                           Z => n8795);
   U4971 : MUX2_X1 port map( A => REGISTERS_77_16_port, B => n2776, S => n1462,
                           Z => n8796);
   U4972 : MUX2_X1 port map( A => REGISTERS_77_15_port, B => n2765, S => n1462,
                           Z => n8797);
   U4973 : MUX2_X1 port map( A => REGISTERS_77_14_port, B => n2754, S => n1462,
                           Z => n8798);
   U4974 : MUX2_X1 port map( A => REGISTERS_77_13_port, B => n2743, S => n1462,
                           Z => n8799);
   U4975 : MUX2_X1 port map( A => REGISTERS_77_12_port, B => n2732, S => n1462,
                           Z => n8800);
   U4976 : MUX2_X1 port map( A => REGISTERS_77_11_port, B => n2721, S => n1462,
                           Z => n8801);
   U4977 : MUX2_X1 port map( A => REGISTERS_77_10_port, B => n2710, S => n1462,
                           Z => n8802);
   U4978 : MUX2_X1 port map( A => REGISTERS_77_9_port, B => n2603, S => n1462, 
                           Z => n8803);
   U4979 : MUX2_X1 port map( A => REGISTERS_77_8_port, B => n2592, S => n1462, 
                           Z => n8804);
   U4980 : MUX2_X1 port map( A => REGISTERS_77_7_port, B => n2581, S => n1463, 
                           Z => n8805);
   U4981 : MUX2_X1 port map( A => REGISTERS_77_6_port, B => n2570, S => n1463, 
                           Z => n8806);
   U4982 : MUX2_X1 port map( A => REGISTERS_77_5_port, B => n2559, S => n1463, 
                           Z => n8807);
   U4983 : MUX2_X1 port map( A => REGISTERS_77_4_port, B => n2548, S => n1463, 
                           Z => n8808);
   U4984 : MUX2_X1 port map( A => REGISTERS_77_3_port, B => n1833, S => n1463, 
                           Z => n8809);
   U4985 : MUX2_X1 port map( A => REGISTERS_77_2_port, B => n1822, S => n1463, 
                           Z => n8810);
   U4986 : MUX2_X1 port map( A => REGISTERS_77_1_port, B => n1811, S => n1463, 
                           Z => n8811);
   U4987 : MUX2_X1 port map( A => REGISTERS_77_0_port, B => n1800, S => n1463, 
                           Z => n8812);
   U4988 : MUX2_X1 port map( A => n10790, B => n2948, S => n1464, Z => 
                           n8749_port);
   U4989 : MUX2_X1 port map( A => n10791, B => n2937, S => n1464, Z => 
                           n8750_port);
   U4990 : MUX2_X1 port map( A => n10792, B => n2926, S => n1464, Z => 
                           n8751_port);
   U4991 : MUX2_X1 port map( A => n10793, B => n2910, S => n1464, Z => 
                           n8752_port);
   U4992 : MUX2_X1 port map( A => n10794, B => n2899, S => n1464, Z => 
                           n8753_port);
   U4993 : MUX2_X1 port map( A => n10795, B => n2887, S => n1464, Z => 
                           n8754_port);
   U4994 : MUX2_X1 port map( A => n10796, B => n2876, S => n1464, Z => 
                           n8755_port);
   U4995 : MUX2_X1 port map( A => n10797, B => n2865, S => n1464, Z => 
                           n8756_port);
   U4996 : MUX2_X1 port map( A => n10798, B => n2854, S => n1464, Z => 
                           n8757_port);
   U4997 : MUX2_X1 port map( A => n10799, B => n2843, S => n1464, Z => 
                           n8758_port);
   U4998 : MUX2_X1 port map( A => n10800, B => n2832, S => n1464, Z => 
                           n8759_port);
   U4999 : MUX2_X1 port map( A => n10801, B => n2821, S => n1464, Z => 
                           n8760_port);
   U5000 : MUX2_X1 port map( A => n10802, B => n2810, S => n1465, Z => 
                           n8761_port);
   U5001 : MUX2_X1 port map( A => n10803, B => n2799, S => n1465, Z => 
                           n8762_port);
   U5002 : MUX2_X1 port map( A => n10804, B => n2788, S => n1465, Z => 
                           n8763_port);
   U5003 : MUX2_X1 port map( A => n10805, B => n2777, S => n1465, Z => 
                           n8764_port);
   U5004 : MUX2_X1 port map( A => n10806, B => n2766, S => n1465, Z => 
                           n8765_port);
   U5005 : MUX2_X1 port map( A => n10807, B => n2755, S => n1465, Z => 
                           n8766_port);
   U5006 : MUX2_X1 port map( A => n10808, B => n2744, S => n1465, Z => 
                           n8767_port);
   U5007 : MUX2_X1 port map( A => n10809, B => n2733, S => n1465, Z => n8768);
   U5008 : MUX2_X1 port map( A => n10810, B => n2722, S => n1465, Z => n8769);
   U5009 : MUX2_X1 port map( A => n10811, B => n2711, S => n1465, Z => n8770);
   U5010 : MUX2_X1 port map( A => n10812, B => n2604, S => n1465, Z => n8771);
   U5011 : MUX2_X1 port map( A => n10813, B => n2593, S => n1465, Z => n8772);
   U5012 : MUX2_X1 port map( A => n10814, B => n2582, S => n1466, Z => n8773);
   U5013 : MUX2_X1 port map( A => n10815, B => n2571, S => n1466, Z => n8774);
   U5014 : MUX2_X1 port map( A => n10816, B => n2560, S => n1466, Z => n8775);
   U5015 : MUX2_X1 port map( A => n10817, B => n2549, S => n1466, Z => n8776);
   U5016 : MUX2_X1 port map( A => n10818, B => n1834, S => n1466, Z => n8777);
   U5017 : MUX2_X1 port map( A => n10819, B => n1823, S => n1466, Z => n8778);
   U5018 : MUX2_X1 port map( A => n10820, B => n1812, S => n1466, Z => n8779);
   U5019 : MUX2_X1 port map( A => n10821, B => n1801, S => n1466, Z => n8780);
   U5020 : MUX2_X1 port map( A => n10758, B => n2948, S => n1467, Z => 
                           n8717_port);
   U5021 : MUX2_X1 port map( A => n10759, B => n2937, S => n1467, Z => 
                           n8718_port);
   U5022 : MUX2_X1 port map( A => n10760, B => n2926, S => n1467, Z => 
                           n8719_port);
   U5023 : MUX2_X1 port map( A => n10761, B => n2910, S => n1467, Z => 
                           n8720_port);
   U5024 : MUX2_X1 port map( A => n10762, B => n2899, S => n1467, Z => 
                           n8721_port);
   U5025 : MUX2_X1 port map( A => n10763, B => n2887, S => n1467, Z => 
                           n8722_port);
   U5026 : MUX2_X1 port map( A => n10764, B => n2876, S => n1467, Z => 
                           n8723_port);
   U5027 : MUX2_X1 port map( A => n10765, B => n2865, S => n1467, Z => 
                           n8724_port);
   U5028 : MUX2_X1 port map( A => n10766, B => n2854, S => n1467, Z => 
                           n8725_port);
   U5029 : MUX2_X1 port map( A => n10767, B => n2843, S => n1467, Z => 
                           n8726_port);
   U5030 : MUX2_X1 port map( A => n10768, B => n2832, S => n1467, Z => 
                           n8727_port);
   U5031 : MUX2_X1 port map( A => n10769, B => n2821, S => n1467, Z => 
                           n8728_port);
   U5032 : MUX2_X1 port map( A => n10770, B => n2810, S => n1468, Z => 
                           n8729_port);
   U5033 : MUX2_X1 port map( A => n10771, B => n2799, S => n1468, Z => 
                           n8730_port);
   U5034 : MUX2_X1 port map( A => n10772, B => n2788, S => n1468, Z => 
                           n8731_port);
   U5035 : MUX2_X1 port map( A => n10773, B => n2777, S => n1468, Z => 
                           n8732_port);
   U5036 : MUX2_X1 port map( A => n10774, B => n2766, S => n1468, Z => 
                           n8733_port);
   U5037 : MUX2_X1 port map( A => n10775, B => n2755, S => n1468, Z => 
                           n8734_port);
   U5038 : MUX2_X1 port map( A => n10776, B => n2744, S => n1468, Z => 
                           n8735_port);
   U5039 : MUX2_X1 port map( A => n10777, B => n2733, S => n1468, Z => 
                           n8736_port);
   U5040 : MUX2_X1 port map( A => n10778, B => n2722, S => n1468, Z => 
                           n8737_port);
   U5041 : MUX2_X1 port map( A => n10779, B => n2711, S => n1468, Z => 
                           n8738_port);
   U5042 : MUX2_X1 port map( A => n10780, B => n2604, S => n1468, Z => 
                           n8739_port);
   U5043 : MUX2_X1 port map( A => n10781, B => n2593, S => n1468, Z => 
                           n8740_port);
   U5044 : MUX2_X1 port map( A => n10782, B => n2582, S => n1469, Z => 
                           n8741_port);
   U5045 : MUX2_X1 port map( A => n10783, B => n2571, S => n1469, Z => 
                           n8742_port);
   U5046 : MUX2_X1 port map( A => n10784, B => n2560, S => n1469, Z => 
                           n8743_port);
   U5047 : MUX2_X1 port map( A => n10785, B => n2549, S => n1469, Z => 
                           n8744_port);
   U5048 : MUX2_X1 port map( A => n10786, B => n1834, S => n1469, Z => 
                           n8745_port);
   U5049 : MUX2_X1 port map( A => n10787, B => n1823, S => n1469, Z => 
                           n8746_port);
   U5050 : MUX2_X1 port map( A => n10788, B => n1812, S => n1469, Z => 
                           n8747_port);
   U5051 : MUX2_X1 port map( A => n10789, B => n1801, S => n1469, Z => 
                           n8748_port);
   U5052 : MUX2_X1 port map( A => n10726, B => n2948, S => n1470, Z => n8685);
   U5053 : MUX2_X1 port map( A => n10727, B => n2937, S => n1470, Z => n8686);
   U5054 : MUX2_X1 port map( A => n10728, B => n2926, S => n1470, Z => n8687);
   U5055 : MUX2_X1 port map( A => n10729, B => n2910, S => n1470, Z => n8688);
   U5056 : MUX2_X1 port map( A => n10730, B => n2899, S => n1470, Z => n8689);
   U5057 : MUX2_X1 port map( A => n10731, B => n2887, S => n1470, Z => n8690);
   U5058 : MUX2_X1 port map( A => n10732, B => n2876, S => n1470, Z => n8691);
   U5059 : MUX2_X1 port map( A => n10733, B => n2865, S => n1470, Z => n8692);
   U5060 : MUX2_X1 port map( A => n10734, B => n2854, S => n1470, Z => n8693);
   U5061 : MUX2_X1 port map( A => n10735, B => n2843, S => n1470, Z => n8694);
   U5062 : MUX2_X1 port map( A => n10736, B => n2832, S => n1470, Z => n8695);
   U5063 : MUX2_X1 port map( A => n10737, B => n2821, S => n1470, Z => n8696);
   U5064 : MUX2_X1 port map( A => n10738, B => n2810, S => n1471, Z => n8697);
   U5065 : MUX2_X1 port map( A => n10739, B => n2799, S => n1471, Z => n8698);
   U5066 : MUX2_X1 port map( A => n10740, B => n2788, S => n1471, Z => n8699);
   U5067 : MUX2_X1 port map( A => n10741, B => n2777, S => n1471, Z => n8700);
   U5068 : MUX2_X1 port map( A => n10742, B => n2766, S => n1471, Z => n8701);
   U5069 : MUX2_X1 port map( A => n10743, B => n2755, S => n1471, Z => 
                           n8702_port);
   U5070 : MUX2_X1 port map( A => n10744, B => n2744, S => n1471, Z => 
                           n8703_port);
   U5071 : MUX2_X1 port map( A => n10745, B => n2733, S => n1471, Z => 
                           n8704_port);
   U5072 : MUX2_X1 port map( A => n10746, B => n2722, S => n1471, Z => 
                           n8705_port);
   U5073 : MUX2_X1 port map( A => n10747, B => n2711, S => n1471, Z => 
                           n8706_port);
   U5074 : MUX2_X1 port map( A => n10748, B => n2604, S => n1471, Z => 
                           n8707_port);
   U5075 : MUX2_X1 port map( A => n10749, B => n2593, S => n1471, Z => 
                           n8708_port);
   U5076 : MUX2_X1 port map( A => n10750, B => n2582, S => n1472, Z => 
                           n8709_port);
   U5077 : MUX2_X1 port map( A => n10751, B => n2571, S => n1472, Z => 
                           n8710_port);
   U5078 : MUX2_X1 port map( A => n10752, B => n2560, S => n1472, Z => 
                           n8711_port);
   U5079 : MUX2_X1 port map( A => n10753, B => n2549, S => n1472, Z => 
                           n8712_port);
   U5080 : MUX2_X1 port map( A => n10754, B => n1834, S => n1472, Z => 
                           n8713_port);
   U5081 : MUX2_X1 port map( A => n10755, B => n1823, S => n1472, Z => 
                           n8714_port);
   U5082 : MUX2_X1 port map( A => n10756, B => n1812, S => n1472, Z => 
                           n8715_port);
   U5083 : MUX2_X1 port map( A => n10757, B => n1801, S => n1472, Z => 
                           n8716_port);
   U5084 : MUX2_X1 port map( A => n10694, B => n2948, S => n1473, Z => n8653);
   U5085 : MUX2_X1 port map( A => n10695, B => n2937, S => n1473, Z => n8654);
   U5086 : MUX2_X1 port map( A => n10696, B => n2926, S => n1473, Z => n8655);
   U5087 : MUX2_X1 port map( A => n10697, B => n2910, S => n1473, Z => n8656);
   U5088 : MUX2_X1 port map( A => n10698, B => n2899, S => n1473, Z => n8657);
   U5089 : MUX2_X1 port map( A => n10699, B => n2887, S => n1473, Z => n8658);
   U5090 : MUX2_X1 port map( A => n10700, B => n2876, S => n1473, Z => n8659);
   U5091 : MUX2_X1 port map( A => n10701, B => n2865, S => n1473, Z => n8660);
   U5092 : MUX2_X1 port map( A => n10702, B => n2854, S => n1473, Z => n8661);
   U5093 : MUX2_X1 port map( A => n10703, B => n2843, S => n1473, Z => n8662);
   U5094 : MUX2_X1 port map( A => n10704, B => n2832, S => n1473, Z => n8663);
   U5095 : MUX2_X1 port map( A => n10705, B => n2821, S => n1473, Z => n8664);
   U5096 : MUX2_X1 port map( A => n10706, B => n2810, S => n1474, Z => n8665);
   U5097 : MUX2_X1 port map( A => n10707, B => n2799, S => n1474, Z => n8666);
   U5098 : MUX2_X1 port map( A => n10708, B => n2788, S => n1474, Z => n8667);
   U5099 : MUX2_X1 port map( A => n10709, B => n2777, S => n1474, Z => n8668);
   U5100 : MUX2_X1 port map( A => n10710, B => n2766, S => n1474, Z => n8669);
   U5101 : MUX2_X1 port map( A => n10711, B => n2755, S => n1474, Z => n8670);
   U5102 : MUX2_X1 port map( A => n10712, B => n2744, S => n1474, Z => n8671);
   U5103 : MUX2_X1 port map( A => n10713, B => n2733, S => n1474, Z => n8672);
   U5104 : MUX2_X1 port map( A => n10714, B => n2722, S => n1474, Z => n8673);
   U5105 : MUX2_X1 port map( A => n10715, B => n2711, S => n1474, Z => n8674);
   U5106 : MUX2_X1 port map( A => n10716, B => n2604, S => n1474, Z => n8675);
   U5107 : MUX2_X1 port map( A => n10717, B => n2593, S => n1474, Z => n8676);
   U5108 : MUX2_X1 port map( A => n10718, B => n2582, S => n1475, Z => n8677);
   U5109 : MUX2_X1 port map( A => n10719, B => n2571, S => n1475, Z => n8678);
   U5110 : MUX2_X1 port map( A => n10720, B => n2560, S => n1475, Z => n8679);
   U5111 : MUX2_X1 port map( A => n10721, B => n2549, S => n1475, Z => n8680);
   U5112 : MUX2_X1 port map( A => n10722, B => n1834, S => n1475, Z => n8681);
   U5113 : MUX2_X1 port map( A => n10723, B => n1823, S => n1475, Z => n8682);
   U5114 : MUX2_X1 port map( A => n10724, B => n1812, S => n1475, Z => n8683);
   U5115 : MUX2_X1 port map( A => n10725, B => n1801, S => n1475, Z => n8684);
   U5116 : MUX2_X1 port map( A => n10662, B => n2948, S => n1476, Z => n8621);
   U5117 : MUX2_X1 port map( A => n10663, B => n2937, S => n1476, Z => n8622);
   U5118 : MUX2_X1 port map( A => n10664, B => n2926, S => n1476, Z => n8623);
   U5119 : MUX2_X1 port map( A => n10665, B => n2910, S => n1476, Z => n8624);
   U5120 : MUX2_X1 port map( A => n10666, B => n2899, S => n1476, Z => n8625);
   U5121 : MUX2_X1 port map( A => n10667, B => n2887, S => n1476, Z => n8626);
   U5122 : MUX2_X1 port map( A => n10668, B => n2876, S => n1476, Z => n8627);
   U5123 : MUX2_X1 port map( A => n10669, B => n2865, S => n1476, Z => n8628);
   U5124 : MUX2_X1 port map( A => n10670, B => n2854, S => n1476, Z => n8629);
   U5125 : MUX2_X1 port map( A => n10671, B => n2843, S => n1476, Z => n8630);
   U5126 : MUX2_X1 port map( A => n10672, B => n2832, S => n1476, Z => n8631);
   U5127 : MUX2_X1 port map( A => n10673, B => n2821, S => n1476, Z => n8632);
   U5128 : MUX2_X1 port map( A => n10674, B => n2810, S => n1477, Z => n8633);
   U5129 : MUX2_X1 port map( A => n10675, B => n2799, S => n1477, Z => n8634);
   U5130 : MUX2_X1 port map( A => n10676, B => n2788, S => n1477, Z => n8635);
   U5131 : MUX2_X1 port map( A => n10677, B => n2777, S => n1477, Z => n8636);
   U5132 : MUX2_X1 port map( A => n10678, B => n2766, S => n1477, Z => n8637);
   U5133 : MUX2_X1 port map( A => n10679, B => n2755, S => n1477, Z => n8638);
   U5134 : MUX2_X1 port map( A => n10680, B => n2744, S => n1477, Z => n8639);
   U5135 : MUX2_X1 port map( A => n10681, B => n2733, S => n1477, Z => n8640);
   U5136 : MUX2_X1 port map( A => n10682, B => n2722, S => n1477, Z => n8641);
   U5137 : MUX2_X1 port map( A => n10683, B => n2711, S => n1477, Z => n8642);
   U5138 : MUX2_X1 port map( A => n10684, B => n2604, S => n1477, Z => n8643);
   U5139 : MUX2_X1 port map( A => n10685, B => n2593, S => n1477, Z => n8644);
   U5140 : MUX2_X1 port map( A => n10686, B => n2582, S => n1478, Z => n8645);
   U5141 : MUX2_X1 port map( A => n10687, B => n2571, S => n1478, Z => n8646);
   U5142 : MUX2_X1 port map( A => n10688, B => n2560, S => n1478, Z => n8647);
   U5143 : MUX2_X1 port map( A => n10689, B => n2549, S => n1478, Z => n8648);
   U5144 : MUX2_X1 port map( A => n10690, B => n1834, S => n1478, Z => n8649);
   U5145 : MUX2_X1 port map( A => n10691, B => n1823, S => n1478, Z => n8650);
   U5146 : MUX2_X1 port map( A => n10692, B => n1812, S => n1478, Z => n8651);
   U5147 : MUX2_X1 port map( A => n10693, B => n1801, S => n1478, Z => n8652);
   U5148 : MUX2_X1 port map( A => n10630, B => n2948, S => n1479, Z => n8589);
   U5149 : MUX2_X1 port map( A => n10631, B => n2937, S => n1479, Z => n8590);
   U5150 : MUX2_X1 port map( A => n10632, B => n2926, S => n1479, Z => n8591);
   U5151 : MUX2_X1 port map( A => n10633, B => n2910, S => n1479, Z => n8592);
   U5152 : MUX2_X1 port map( A => n10634, B => n2899, S => n1479, Z => n8593);
   U5153 : MUX2_X1 port map( A => n10635, B => n2887, S => n1479, Z => n8594);
   U5154 : MUX2_X1 port map( A => n10636, B => n2876, S => n1479, Z => n8595);
   U5155 : MUX2_X1 port map( A => n10637, B => n2865, S => n1479, Z => n8596);
   U5156 : MUX2_X1 port map( A => n10638, B => n2854, S => n1479, Z => n8597);
   U5157 : MUX2_X1 port map( A => n10639, B => n2843, S => n1479, Z => n8598);
   U5158 : MUX2_X1 port map( A => n10640, B => n2832, S => n1479, Z => n8599);
   U5159 : MUX2_X1 port map( A => n10641, B => n2821, S => n1479, Z => n8600);
   U5160 : MUX2_X1 port map( A => n10642, B => n2810, S => n1480, Z => n8601);
   U5161 : MUX2_X1 port map( A => n10643, B => n2799, S => n1480, Z => n8602);
   U5162 : MUX2_X1 port map( A => n10644, B => n2788, S => n1480, Z => n8603);
   U5163 : MUX2_X1 port map( A => n10645, B => n2777, S => n1480, Z => n8604);
   U5164 : MUX2_X1 port map( A => n10646, B => n2766, S => n1480, Z => n8605);
   U5165 : MUX2_X1 port map( A => n10647, B => n2755, S => n1480, Z => n8606);
   U5166 : MUX2_X1 port map( A => n10648, B => n2744, S => n1480, Z => n8607);
   U5167 : MUX2_X1 port map( A => n10649, B => n2733, S => n1480, Z => n8608);
   U5168 : MUX2_X1 port map( A => n10650, B => n2722, S => n1480, Z => n8609);
   U5169 : MUX2_X1 port map( A => n10651, B => n2711, S => n1480, Z => n8610);
   U5170 : MUX2_X1 port map( A => n10652, B => n2604, S => n1480, Z => n8611);
   U5171 : MUX2_X1 port map( A => n10653, B => n2593, S => n1480, Z => n8612);
   U5172 : MUX2_X1 port map( A => n10654, B => n2582, S => n1481, Z => n8613);
   U5173 : MUX2_X1 port map( A => n10655, B => n2571, S => n1481, Z => n8614);
   U5174 : MUX2_X1 port map( A => n10656, B => n2560, S => n1481, Z => n8615);
   U5175 : MUX2_X1 port map( A => n10657, B => n2549, S => n1481, Z => n8616);
   U5176 : MUX2_X1 port map( A => n10658, B => n1834, S => n1481, Z => n8617);
   U5177 : MUX2_X1 port map( A => n10659, B => n1823, S => n1481, Z => n8618);
   U5178 : MUX2_X1 port map( A => n10660, B => n1812, S => n1481, Z => n8619);
   U5179 : MUX2_X1 port map( A => n10661, B => n1801, S => n1481, Z => n8620);
   U5180 : MUX2_X1 port map( A => n10598, B => n2948, S => n1482, Z => n8557);
   U5181 : MUX2_X1 port map( A => n10599, B => n2937, S => n1482, Z => n8558);
   U5182 : MUX2_X1 port map( A => n10600, B => n2926, S => n1482, Z => 
                           n8559_port);
   U5183 : MUX2_X1 port map( A => n10601, B => n2910, S => n1482, Z => n8560);
   U5184 : MUX2_X1 port map( A => n10602, B => n2899, S => n1482, Z => 
                           n8561_port);
   U5185 : MUX2_X1 port map( A => n10603, B => n2887, S => n1482, Z => 
                           n8562_port);
   U5186 : MUX2_X1 port map( A => n10604, B => n2876, S => n1482, Z => 
                           n8563_port);
   U5187 : MUX2_X1 port map( A => n10605, B => n2865, S => n1482, Z => 
                           n8564_port);
   U5188 : MUX2_X1 port map( A => n10606, B => n2854, S => n1482, Z => 
                           n8565_port);
   U5189 : MUX2_X1 port map( A => n10607, B => n2843, S => n1482, Z => 
                           n8566_port);
   U5190 : MUX2_X1 port map( A => n10608, B => n2832, S => n1482, Z => 
                           n8567_port);
   U5191 : MUX2_X1 port map( A => n10609, B => n2821, S => n1482, Z => n8568);
   U5192 : MUX2_X1 port map( A => n10610, B => n2810, S => n1483, Z => n8569);
   U5193 : MUX2_X1 port map( A => n10611, B => n2799, S => n1483, Z => n8570);
   U5194 : MUX2_X1 port map( A => n10612, B => n2788, S => n1483, Z => 
                           n8571_port);
   U5195 : MUX2_X1 port map( A => n10613, B => n2777, S => n1483, Z => 
                           n8572_port);
   U5196 : MUX2_X1 port map( A => n10614, B => n2766, S => n1483, Z => 
                           n8573_port);
   U5197 : MUX2_X1 port map( A => n10615, B => n2755, S => n1483, Z => 
                           n8574_port);
   U5198 : MUX2_X1 port map( A => n10616, B => n2744, S => n1483, Z => n8575);
   U5199 : MUX2_X1 port map( A => n10617, B => n2733, S => n1483, Z => n8576);
   U5200 : MUX2_X1 port map( A => n10618, B => n2722, S => n1483, Z => n8577);
   U5201 : MUX2_X1 port map( A => n10619, B => n2711, S => n1483, Z => n8578);
   U5202 : MUX2_X1 port map( A => n10620, B => n2604, S => n1483, Z => n8579);
   U5203 : MUX2_X1 port map( A => n10621, B => n2593, S => n1483, Z => n8580);
   U5204 : MUX2_X1 port map( A => n10622, B => n2582, S => n1484, Z => n8581);
   U5205 : MUX2_X1 port map( A => n10623, B => n2571, S => n1484, Z => n8582);
   U5206 : MUX2_X1 port map( A => n10624, B => n2560, S => n1484, Z => n8583);
   U5207 : MUX2_X1 port map( A => n10625, B => n2549, S => n1484, Z => n8584);
   U5208 : MUX2_X1 port map( A => n10626, B => n1834, S => n1484, Z => n8585);
   U5209 : MUX2_X1 port map( A => n10627, B => n1823, S => n1484, Z => n8586);
   U5210 : MUX2_X1 port map( A => n10628, B => n1812, S => n1484, Z => n8587);
   U5211 : MUX2_X1 port map( A => n10629, B => n1801, S => n1484, Z => n8588);
   U5212 : MUX2_X1 port map( A => n10566, B => n2948, S => n1485, Z => n8525);
   U5213 : MUX2_X1 port map( A => n10567, B => n2937, S => n1485, Z => n8526);
   U5214 : MUX2_X1 port map( A => n10568, B => n2926, S => n1485, Z => n8527);
   U5215 : MUX2_X1 port map( A => n10569, B => n2910, S => n1485, Z => n8528);
   U5216 : MUX2_X1 port map( A => n10570, B => n2899, S => n1485, Z => n8529);
   U5217 : MUX2_X1 port map( A => n10571, B => n2887, S => n1485, Z => n8530);
   U5218 : MUX2_X1 port map( A => n10572, B => n2876, S => n1485, Z => n8531);
   U5219 : MUX2_X1 port map( A => n10573, B => n2865, S => n1485, Z => n8532);
   U5220 : MUX2_X1 port map( A => n10574, B => n2854, S => n1485, Z => n8533);
   U5221 : MUX2_X1 port map( A => n10575, B => n2843, S => n1485, Z => n8534);
   U5222 : MUX2_X1 port map( A => n10576, B => n2832, S => n1485, Z => n8535);
   U5223 : MUX2_X1 port map( A => n10577, B => n2821, S => n1485, Z => n8536);
   U5224 : MUX2_X1 port map( A => n10578, B => n2810, S => n1486, Z => n8537);
   U5225 : MUX2_X1 port map( A => n10579, B => n2799, S => n1486, Z => n8538);
   U5226 : MUX2_X1 port map( A => n10580, B => n2788, S => n1486, Z => n8539);
   U5227 : MUX2_X1 port map( A => n10581, B => n2777, S => n1486, Z => n8540);
   U5228 : MUX2_X1 port map( A => n10582, B => n2766, S => n1486, Z => n8541);
   U5229 : MUX2_X1 port map( A => n10583, B => n2755, S => n1486, Z => n8542);
   U5230 : MUX2_X1 port map( A => n10584, B => n2744, S => n1486, Z => n8543);
   U5231 : MUX2_X1 port map( A => n10585, B => n2733, S => n1486, Z => n8544);
   U5232 : MUX2_X1 port map( A => n10586, B => n2722, S => n1486, Z => n8545);
   U5233 : MUX2_X1 port map( A => n10587, B => n2711, S => n1486, Z => n8546);
   U5234 : MUX2_X1 port map( A => n10588, B => n2604, S => n1486, Z => n8547);
   U5235 : MUX2_X1 port map( A => n10589, B => n2593, S => n1486, Z => n8548);
   U5236 : MUX2_X1 port map( A => n10590, B => n2582, S => n1487, Z => n8549);
   U5237 : MUX2_X1 port map( A => n10591, B => n2571, S => n1487, Z => n8550);
   U5238 : MUX2_X1 port map( A => n10592, B => n2560, S => n1487, Z => n8551);
   U5239 : MUX2_X1 port map( A => n10593, B => n2549, S => n1487, Z => n8552);
   U5240 : MUX2_X1 port map( A => n10594, B => n1834, S => n1487, Z => n8553);
   U5241 : MUX2_X1 port map( A => n10595, B => n1823, S => n1487, Z => n8554);
   U5242 : MUX2_X1 port map( A => n10596, B => n1812, S => n1487, Z => n8555);
   U5243 : MUX2_X1 port map( A => n10597, B => n1801, S => n1487, Z => n8556);
   U5244 : MUX2_X1 port map( A => n10534, B => n2948, S => n1488, Z => n8493);
   U5245 : MUX2_X1 port map( A => n10535, B => n2937, S => n1488, Z => n8494);
   U5246 : MUX2_X1 port map( A => n10536, B => n2926, S => n1488, Z => n8495);
   U5247 : MUX2_X1 port map( A => n10537, B => n2910, S => n1488, Z => n8496);
   U5248 : MUX2_X1 port map( A => n10538, B => n2899, S => n1488, Z => n8497);
   U5249 : MUX2_X1 port map( A => n10539, B => n2887, S => n1488, Z => n8498);
   U5250 : MUX2_X1 port map( A => n10540, B => n2876, S => n1488, Z => n8499);
   U5251 : MUX2_X1 port map( A => n10541, B => n2865, S => n1488, Z => n8500);
   U5252 : MUX2_X1 port map( A => n10542, B => n2854, S => n1488, Z => n8501);
   U5253 : MUX2_X1 port map( A => n10543, B => n2843, S => n1488, Z => n8502);
   U5254 : MUX2_X1 port map( A => n10544, B => n2832, S => n1488, Z => n8503);
   U5255 : MUX2_X1 port map( A => n10545, B => n2821, S => n1488, Z => n8504);
   U5256 : MUX2_X1 port map( A => n10546, B => n2810, S => n1489, Z => n8505);
   U5257 : MUX2_X1 port map( A => n10547, B => n2799, S => n1489, Z => n8506);
   U5258 : MUX2_X1 port map( A => n10548, B => n2788, S => n1489, Z => n8507);
   U5259 : MUX2_X1 port map( A => n10549, B => n2777, S => n1489, Z => n8508);
   U5260 : MUX2_X1 port map( A => n10550, B => n2766, S => n1489, Z => n8509);
   U5261 : MUX2_X1 port map( A => n10551, B => n2755, S => n1489, Z => n8510);
   U5262 : MUX2_X1 port map( A => n10552, B => n2744, S => n1489, Z => n8511);
   U5263 : MUX2_X1 port map( A => n10553, B => n2733, S => n1489, Z => n8512);
   U5264 : MUX2_X1 port map( A => n10554, B => n2722, S => n1489, Z => n8513);
   U5265 : MUX2_X1 port map( A => n10555, B => n2711, S => n1489, Z => n8514);
   U5266 : MUX2_X1 port map( A => n10556, B => n2604, S => n1489, Z => n8515);
   U5267 : MUX2_X1 port map( A => n10557, B => n2593, S => n1489, Z => n8516);
   U5268 : MUX2_X1 port map( A => n10558, B => n2582, S => n1490, Z => n8517);
   U5269 : MUX2_X1 port map( A => n10559, B => n2571, S => n1490, Z => n8518);
   U5270 : MUX2_X1 port map( A => n10560, B => n2560, S => n1490, Z => n8519);
   U5271 : MUX2_X1 port map( A => n10561, B => n2549, S => n1490, Z => n8520);
   U5272 : MUX2_X1 port map( A => n10562, B => n1834, S => n1490, Z => n8521);
   U5273 : MUX2_X1 port map( A => n10563, B => n1823, S => n1490, Z => n8522);
   U5274 : MUX2_X1 port map( A => n10564, B => n1812, S => n1490, Z => n8523);
   U5275 : MUX2_X1 port map( A => n10565, B => n1801, S => n1490, Z => n8524);
   U5276 : MUX2_X1 port map( A => n10502, B => n2948, S => n1491, Z => n8461);
   U5277 : MUX2_X1 port map( A => n10503, B => n2937, S => n1491, Z => n8462);
   U5278 : MUX2_X1 port map( A => n10504, B => n2926, S => n1491, Z => n8463);
   U5279 : MUX2_X1 port map( A => n10505, B => n2910, S => n1491, Z => n8464);
   U5280 : MUX2_X1 port map( A => n10506, B => n2899, S => n1491, Z => n8465);
   U5281 : MUX2_X1 port map( A => n10507, B => n2887, S => n1491, Z => n8466);
   U5282 : MUX2_X1 port map( A => n10508, B => n2876, S => n1491, Z => n8467);
   U5283 : MUX2_X1 port map( A => n10509, B => n2865, S => n1491, Z => n8468);
   U5284 : MUX2_X1 port map( A => n10510, B => n2854, S => n1491, Z => n8469);
   U5285 : MUX2_X1 port map( A => n10511, B => n2843, S => n1491, Z => n8470);
   U5286 : MUX2_X1 port map( A => n10512, B => n2832, S => n1491, Z => n8471);
   U5287 : MUX2_X1 port map( A => n10513, B => n2821, S => n1491, Z => n8472);
   U5288 : MUX2_X1 port map( A => n10514, B => n2810, S => n1492, Z => n8473);
   U5289 : MUX2_X1 port map( A => n10515, B => n2799, S => n1492, Z => n8474);
   U5290 : MUX2_X1 port map( A => n10516, B => n2788, S => n1492, Z => n8475);
   U5291 : MUX2_X1 port map( A => n10517, B => n2777, S => n1492, Z => n8476);
   U5292 : MUX2_X1 port map( A => n10518, B => n2766, S => n1492, Z => n8477);
   U5293 : MUX2_X1 port map( A => n10519, B => n2755, S => n1492, Z => n8478);
   U5294 : MUX2_X1 port map( A => n10520, B => n2744, S => n1492, Z => n8479);
   U5295 : MUX2_X1 port map( A => n10521, B => n2733, S => n1492, Z => n8480);
   U5296 : MUX2_X1 port map( A => n10522, B => n2722, S => n1492, Z => n8481);
   U5297 : MUX2_X1 port map( A => n10523, B => n2711, S => n1492, Z => n8482);
   U5298 : MUX2_X1 port map( A => n10524, B => n2604, S => n1492, Z => n8483);
   U5299 : MUX2_X1 port map( A => n10525, B => n2593, S => n1492, Z => n8484);
   U5300 : MUX2_X1 port map( A => n10526, B => n2582, S => n1493, Z => n8485);
   U5301 : MUX2_X1 port map( A => n10527, B => n2571, S => n1493, Z => n8486);
   U5302 : MUX2_X1 port map( A => n10528, B => n2560, S => n1493, Z => n8487);
   U5303 : MUX2_X1 port map( A => n10529, B => n2549, S => n1493, Z => n8488);
   U5304 : MUX2_X1 port map( A => n10530, B => n1834, S => n1493, Z => n8489);
   U5305 : MUX2_X1 port map( A => n10531, B => n1823, S => n1493, Z => n8490);
   U5306 : MUX2_X1 port map( A => n10532, B => n1812, S => n1493, Z => n8491);
   U5307 : MUX2_X1 port map( A => n10533, B => n1801, S => n1493, Z => n8492);
   U5308 : MUX2_X1 port map( A => n10470, B => n2948, S => n1494, Z => 
                           n8429_port);
   U5309 : MUX2_X1 port map( A => n10471, B => n2937, S => n1494, Z => 
                           n8430_port);
   U5310 : MUX2_X1 port map( A => n10472, B => n2926, S => n1494, Z => n8431);
   U5311 : MUX2_X1 port map( A => n10473, B => n2910, S => n1494, Z => n8432);
   U5312 : MUX2_X1 port map( A => n10474, B => n2899, S => n1494, Z => n8433);
   U5313 : MUX2_X1 port map( A => n10475, B => n2887, S => n1494, Z => n8434);
   U5314 : MUX2_X1 port map( A => n10476, B => n2876, S => n1494, Z => n8435);
   U5315 : MUX2_X1 port map( A => n10477, B => n2865, S => n1494, Z => n8436);
   U5316 : MUX2_X1 port map( A => n10478, B => n2854, S => n1494, Z => n8437);
   U5317 : MUX2_X1 port map( A => n10479, B => n2843, S => n1494, Z => n8438);
   U5318 : MUX2_X1 port map( A => n10480, B => n2832, S => n1494, Z => n8439);
   U5319 : MUX2_X1 port map( A => n10481, B => n2821, S => n1494, Z => n8440);
   U5320 : MUX2_X1 port map( A => n10482, B => n2810, S => n1495, Z => n8441);
   U5321 : MUX2_X1 port map( A => n10483, B => n2799, S => n1495, Z => n8442);
   U5322 : MUX2_X1 port map( A => n10484, B => n2788, S => n1495, Z => n8443);
   U5323 : MUX2_X1 port map( A => n10485, B => n2777, S => n1495, Z => n8444);
   U5324 : MUX2_X1 port map( A => n10486, B => n2766, S => n1495, Z => n8445);
   U5325 : MUX2_X1 port map( A => n10487, B => n2755, S => n1495, Z => n8446);
   U5326 : MUX2_X1 port map( A => n10488, B => n2744, S => n1495, Z => n8447);
   U5327 : MUX2_X1 port map( A => n10489, B => n2733, S => n1495, Z => n8448);
   U5328 : MUX2_X1 port map( A => n10490, B => n2722, S => n1495, Z => n8449);
   U5329 : MUX2_X1 port map( A => n10491, B => n2711, S => n1495, Z => n8450);
   U5330 : MUX2_X1 port map( A => n10492, B => n2604, S => n1495, Z => n8451);
   U5331 : MUX2_X1 port map( A => n10493, B => n2593, S => n1495, Z => n8452);
   U5332 : MUX2_X1 port map( A => n10494, B => n2582, S => n1496, Z => n8453);
   U5333 : MUX2_X1 port map( A => n10495, B => n2571, S => n1496, Z => n8454);
   U5334 : MUX2_X1 port map( A => n10496, B => n2560, S => n1496, Z => n8455);
   U5335 : MUX2_X1 port map( A => n10497, B => n2549, S => n1496, Z => n8456);
   U5336 : MUX2_X1 port map( A => n10498, B => n1834, S => n1496, Z => n8457);
   U5337 : MUX2_X1 port map( A => n10499, B => n1823, S => n1496, Z => n8458);
   U5338 : MUX2_X1 port map( A => n10500, B => n1812, S => n1496, Z => n8459);
   U5339 : MUX2_X1 port map( A => n10501, B => n1801, S => n1496, Z => n8460);
   U5340 : MUX2_X1 port map( A => n10438, B => n2949, S => n1497, Z => n8397);
   U5341 : MUX2_X1 port map( A => n10439, B => n2938, S => n1497, Z => n8398);
   U5342 : MUX2_X1 port map( A => n10440, B => n2927, S => n1497, Z => n8399);
   U5343 : MUX2_X1 port map( A => n10441, B => n2911, S => n1497, Z => n8400);
   U5344 : MUX2_X1 port map( A => n10442, B => n2900, S => n1497, Z => n8401);
   U5345 : MUX2_X1 port map( A => n10443, B => n2888, S => n1497, Z => n8402);
   U5346 : MUX2_X1 port map( A => n10444, B => n2877, S => n1497, Z => n8403);
   U5347 : MUX2_X1 port map( A => n10445, B => n2866, S => n1497, Z => n8404);
   U5348 : MUX2_X1 port map( A => n10446, B => n2855, S => n1497, Z => n8405);
   U5349 : MUX2_X1 port map( A => n10447, B => n2844, S => n1497, Z => n8406);
   U5350 : MUX2_X1 port map( A => n10448, B => n2833, S => n1497, Z => n8407);
   U5351 : MUX2_X1 port map( A => n10449, B => n2822, S => n1497, Z => n8408);
   U5352 : MUX2_X1 port map( A => n10450, B => n2811, S => n1498, Z => n8409);
   U5353 : MUX2_X1 port map( A => n10451, B => n2800, S => n1498, Z => n8410);
   U5354 : MUX2_X1 port map( A => n10452, B => n2789, S => n1498, Z => n8411);
   U5355 : MUX2_X1 port map( A => n10453, B => n2778, S => n1498, Z => n8412);
   U5356 : MUX2_X1 port map( A => n10454, B => n2767, S => n1498, Z => n8413);
   U5357 : MUX2_X1 port map( A => n10455, B => n2756, S => n1498, Z => n8414);
   U5358 : MUX2_X1 port map( A => n10456, B => n2745, S => n1498, Z => 
                           n8415_port);
   U5359 : MUX2_X1 port map( A => n10457, B => n2734, S => n1498, Z => n8416);
   U5360 : MUX2_X1 port map( A => n10458, B => n2723, S => n1498, Z => 
                           n8417_port);
   U5361 : MUX2_X1 port map( A => n10459, B => n2712, S => n1498, Z => 
                           n8418_port);
   U5362 : MUX2_X1 port map( A => n10460, B => n2605, S => n1498, Z => 
                           n8419_port);
   U5363 : MUX2_X1 port map( A => n10461, B => n2594, S => n1498, Z => 
                           n8420_port);
   U5364 : MUX2_X1 port map( A => n10462, B => n2583, S => n1499, Z => 
                           n8421_port);
   U5365 : MUX2_X1 port map( A => n10463, B => n2572, S => n1499, Z => 
                           n8422_port);
   U5366 : MUX2_X1 port map( A => n10464, B => n2561, S => n1499, Z => 
                           n8423_port);
   U5367 : MUX2_X1 port map( A => n10465, B => n2550, S => n1499, Z => n8424);
   U5368 : MUX2_X1 port map( A => n10466, B => n1835, S => n1499, Z => n8425);
   U5369 : MUX2_X1 port map( A => n10467, B => n1824, S => n1499, Z => n8426);
   U5370 : MUX2_X1 port map( A => n10468, B => n1813, S => n1499, Z => 
                           n8427_port);
   U5371 : MUX2_X1 port map( A => n10469, B => n1802, S => n1499, Z => 
                           n8428_port);
   U5372 : MUX2_X1 port map( A => n10406, B => n2949, S => n1500, Z => n8365);
   U5373 : MUX2_X1 port map( A => n10407, B => n2938, S => n1500, Z => n8366);
   U5374 : MUX2_X1 port map( A => n10408, B => n2927, S => n1500, Z => n8367);
   U5375 : MUX2_X1 port map( A => n10409, B => n2911, S => n1500, Z => n8368);
   U5376 : MUX2_X1 port map( A => n10410, B => n2900, S => n1500, Z => n8369);
   U5377 : MUX2_X1 port map( A => n10411, B => n2888, S => n1500, Z => n8370);
   U5378 : MUX2_X1 port map( A => n10412, B => n2877, S => n1500, Z => n8371);
   U5379 : MUX2_X1 port map( A => n10413, B => n2866, S => n1500, Z => n8372);
   U5380 : MUX2_X1 port map( A => n10414, B => n2855, S => n1500, Z => n8373);
   U5381 : MUX2_X1 port map( A => n10415, B => n2844, S => n1500, Z => n8374);
   U5382 : MUX2_X1 port map( A => n10416, B => n2833, S => n1500, Z => n8375);
   U5383 : MUX2_X1 port map( A => n10417, B => n2822, S => n1500, Z => n8376);
   U5384 : MUX2_X1 port map( A => n10418, B => n2811, S => n1501, Z => n8377);
   U5385 : MUX2_X1 port map( A => n10419, B => n2800, S => n1501, Z => n8378);
   U5386 : MUX2_X1 port map( A => n10420, B => n2789, S => n1501, Z => n8379);
   U5387 : MUX2_X1 port map( A => n10421, B => n2778, S => n1501, Z => n8380);
   U5388 : MUX2_X1 port map( A => n10422, B => n2767, S => n1501, Z => n8381);
   U5389 : MUX2_X1 port map( A => n10423, B => n2756, S => n1501, Z => n8382);
   U5390 : MUX2_X1 port map( A => n10424, B => n2745, S => n1501, Z => n8383);
   U5391 : MUX2_X1 port map( A => n10425, B => n2734, S => n1501, Z => n8384);
   U5392 : MUX2_X1 port map( A => n10426, B => n2723, S => n1501, Z => n8385);
   U5393 : MUX2_X1 port map( A => n10427, B => n2712, S => n1501, Z => n8386);
   U5394 : MUX2_X1 port map( A => n10428, B => n2605, S => n1501, Z => n8387);
   U5395 : MUX2_X1 port map( A => n10429, B => n2594, S => n1501, Z => n8388);
   U5396 : MUX2_X1 port map( A => n10430, B => n2583, S => n1502, Z => n8389);
   U5397 : MUX2_X1 port map( A => n10431, B => n2572, S => n1502, Z => n8390);
   U5398 : MUX2_X1 port map( A => n10432, B => n2561, S => n1502, Z => n8391);
   U5399 : MUX2_X1 port map( A => n10433, B => n2550, S => n1502, Z => n8392);
   U5400 : MUX2_X1 port map( A => n10434, B => n1835, S => n1502, Z => n8393);
   U5401 : MUX2_X1 port map( A => n10435, B => n1824, S => n1502, Z => n8394);
   U5402 : MUX2_X1 port map( A => n10436, B => n1813, S => n1502, Z => n8395);
   U5403 : MUX2_X1 port map( A => n10437, B => n1802, S => n1502, Z => n8396);
   U5404 : MUX2_X1 port map( A => n10374, B => n2949, S => n1503, Z => n8333);
   U5405 : MUX2_X1 port map( A => n10375, B => n2938, S => n1503, Z => n8334);
   U5406 : MUX2_X1 port map( A => n10376, B => n2927, S => n1503, Z => n8335);
   U5407 : MUX2_X1 port map( A => n10377, B => n2911, S => n1503, Z => n8336);
   U5408 : MUX2_X1 port map( A => n10378, B => n2900, S => n1503, Z => n8337);
   U5409 : MUX2_X1 port map( A => n10379, B => n2888, S => n1503, Z => n8338);
   U5410 : MUX2_X1 port map( A => n10380, B => n2877, S => n1503, Z => n8339);
   U5411 : MUX2_X1 port map( A => n10381, B => n2866, S => n1503, Z => n8340);
   U5412 : MUX2_X1 port map( A => n10382, B => n2855, S => n1503, Z => n8341);
   U5413 : MUX2_X1 port map( A => n10383, B => n2844, S => n1503, Z => n8342);
   U5414 : MUX2_X1 port map( A => n10384, B => n2833, S => n1503, Z => n8343);
   U5415 : MUX2_X1 port map( A => n10385, B => n2822, S => n1503, Z => n8344);
   U5416 : MUX2_X1 port map( A => n10386, B => n2811, S => n1504, Z => n8345);
   U5417 : MUX2_X1 port map( A => n10387, B => n2800, S => n1504, Z => n8346);
   U5418 : MUX2_X1 port map( A => n10388, B => n2789, S => n1504, Z => n8347);
   U5419 : MUX2_X1 port map( A => n10389, B => n2778, S => n1504, Z => n8348);
   U5420 : MUX2_X1 port map( A => n10390, B => n2767, S => n1504, Z => n8349);
   U5421 : MUX2_X1 port map( A => n10391, B => n2756, S => n1504, Z => n8350);
   U5422 : MUX2_X1 port map( A => n10392, B => n2745, S => n1504, Z => n8351);
   U5423 : MUX2_X1 port map( A => n10393, B => n2734, S => n1504, Z => n8352);
   U5424 : MUX2_X1 port map( A => n10394, B => n2723, S => n1504, Z => n8353);
   U5425 : MUX2_X1 port map( A => n10395, B => n2712, S => n1504, Z => n8354);
   U5426 : MUX2_X1 port map( A => n10396, B => n2605, S => n1504, Z => n8355);
   U5427 : MUX2_X1 port map( A => n10397, B => n2594, S => n1504, Z => n8356);
   U5428 : MUX2_X1 port map( A => n10398, B => n2583, S => n1505, Z => n8357);
   U5429 : MUX2_X1 port map( A => n10399, B => n2572, S => n1505, Z => n8358);
   U5430 : MUX2_X1 port map( A => n10400, B => n2561, S => n1505, Z => n8359);
   U5431 : MUX2_X1 port map( A => n10401, B => n2550, S => n1505, Z => n8360);
   U5432 : MUX2_X1 port map( A => n10402, B => n1835, S => n1505, Z => n8361);
   U5433 : MUX2_X1 port map( A => n10403, B => n1824, S => n1505, Z => n8362);
   U5434 : MUX2_X1 port map( A => n10404, B => n1813, S => n1505, Z => n8363);
   U5435 : MUX2_X1 port map( A => n10405, B => n1802, S => n1505, Z => n8364);
   U5436 : MUX2_X1 port map( A => n10342, B => n2949, S => n1506, Z => n8301);
   U5437 : MUX2_X1 port map( A => n10343, B => n2938, S => n1506, Z => n8302);
   U5438 : MUX2_X1 port map( A => n10344, B => n2927, S => n1506, Z => n8303);
   U5439 : MUX2_X1 port map( A => n10345, B => n2911, S => n1506, Z => n8304);
   U5440 : MUX2_X1 port map( A => n10346, B => n2900, S => n1506, Z => n8305);
   U5441 : MUX2_X1 port map( A => n10347, B => n2888, S => n1506, Z => n8306);
   U5442 : MUX2_X1 port map( A => n10348, B => n2877, S => n1506, Z => n8307);
   U5443 : MUX2_X1 port map( A => n10349, B => n2866, S => n1506, Z => n8308);
   U5444 : MUX2_X1 port map( A => n10350, B => n2855, S => n1506, Z => n8309);
   U5445 : MUX2_X1 port map( A => n10351, B => n2844, S => n1506, Z => n8310);
   U5446 : MUX2_X1 port map( A => n10352, B => n2833, S => n1506, Z => n8311);
   U5447 : MUX2_X1 port map( A => n10353, B => n2822, S => n1506, Z => n8312);
   U5448 : MUX2_X1 port map( A => n10354, B => n2811, S => n1507, Z => n8313);
   U5449 : MUX2_X1 port map( A => n10355, B => n2800, S => n1507, Z => n8314);
   U5450 : MUX2_X1 port map( A => n10356, B => n2789, S => n1507, Z => n8315);
   U5451 : MUX2_X1 port map( A => n10357, B => n2778, S => n1507, Z => n8316);
   U5452 : MUX2_X1 port map( A => n10358, B => n2767, S => n1507, Z => n8317);
   U5453 : MUX2_X1 port map( A => n10359, B => n2756, S => n1507, Z => n8318);
   U5454 : MUX2_X1 port map( A => n10360, B => n2745, S => n1507, Z => n8319);
   U5455 : MUX2_X1 port map( A => n10361, B => n2734, S => n1507, Z => n8320);
   U5456 : MUX2_X1 port map( A => n10362, B => n2723, S => n1507, Z => n8321);
   U5457 : MUX2_X1 port map( A => n10363, B => n2712, S => n1507, Z => n8322);
   U5458 : MUX2_X1 port map( A => n10364, B => n2605, S => n1507, Z => n8323);
   U5459 : MUX2_X1 port map( A => n10365, B => n2594, S => n1507, Z => n8324);
   U5460 : MUX2_X1 port map( A => n10366, B => n2583, S => n1508, Z => n8325);
   U5461 : MUX2_X1 port map( A => n10367, B => n2572, S => n1508, Z => n8326);
   U5462 : MUX2_X1 port map( A => n10368, B => n2561, S => n1508, Z => n8327);
   U5463 : MUX2_X1 port map( A => n10369, B => n2550, S => n1508, Z => n8328);
   U5464 : MUX2_X1 port map( A => n10370, B => n1835, S => n1508, Z => n8329);
   U5465 : MUX2_X1 port map( A => n10371, B => n1824, S => n1508, Z => n8330);
   U5466 : MUX2_X1 port map( A => n10372, B => n1813, S => n1508, Z => n8331);
   U5467 : MUX2_X1 port map( A => n10373, B => n1802, S => n1508, Z => n8332);
   U5468 : MUX2_X1 port map( A => n10310, B => n2949, S => n1509, Z => n8269);
   U5469 : MUX2_X1 port map( A => n10311, B => n2938, S => n1509, Z => n8270);
   U5470 : MUX2_X1 port map( A => n10312, B => n2927, S => n1509, Z => n8271);
   U5471 : MUX2_X1 port map( A => n10313, B => n2911, S => n1509, Z => n8272);
   U5472 : MUX2_X1 port map( A => n10314, B => n2900, S => n1509, Z => n8273);
   U5473 : MUX2_X1 port map( A => n10315, B => n2888, S => n1509, Z => n8274);
   U5474 : MUX2_X1 port map( A => n10316, B => n2877, S => n1509, Z => n8275);
   U5475 : MUX2_X1 port map( A => n10317, B => n2866, S => n1509, Z => n8276);
   U5476 : MUX2_X1 port map( A => n10318, B => n2855, S => n1509, Z => n8277);
   U5477 : MUX2_X1 port map( A => n10319, B => n2844, S => n1509, Z => n8278);
   U5478 : MUX2_X1 port map( A => n10320, B => n2833, S => n1509, Z => n8279);
   U5479 : MUX2_X1 port map( A => n10321, B => n2822, S => n1509, Z => n8280);
   U5480 : MUX2_X1 port map( A => n10322, B => n2811, S => n1510, Z => n8281);
   U5481 : MUX2_X1 port map( A => n10323, B => n2800, S => n1510, Z => n8282);
   U5482 : MUX2_X1 port map( A => n10324, B => n2789, S => n1510, Z => n8283);
   U5483 : MUX2_X1 port map( A => n10325, B => n2778, S => n1510, Z => n8284);
   U5484 : MUX2_X1 port map( A => n10326, B => n2767, S => n1510, Z => n8285);
   U5485 : MUX2_X1 port map( A => n10327, B => n2756, S => n1510, Z => n8286);
   U5486 : MUX2_X1 port map( A => n10328, B => n2745, S => n1510, Z => n8287);
   U5487 : MUX2_X1 port map( A => n10329, B => n2734, S => n1510, Z => n8288);
   U5488 : MUX2_X1 port map( A => n10330, B => n2723, S => n1510, Z => n8289);
   U5489 : MUX2_X1 port map( A => n10331, B => n2712, S => n1510, Z => n8290);
   U5490 : MUX2_X1 port map( A => n10332, B => n2605, S => n1510, Z => n8291);
   U5491 : MUX2_X1 port map( A => n10333, B => n2594, S => n1510, Z => n8292);
   U5492 : MUX2_X1 port map( A => n10334, B => n2583, S => n1511, Z => n8293);
   U5493 : MUX2_X1 port map( A => n10335, B => n2572, S => n1511, Z => n8294);
   U5494 : MUX2_X1 port map( A => n10336, B => n2561, S => n1511, Z => n8295);
   U5495 : MUX2_X1 port map( A => n10337, B => n2550, S => n1511, Z => n8296);
   U5496 : MUX2_X1 port map( A => n10338, B => n1835, S => n1511, Z => n8297);
   U5497 : MUX2_X1 port map( A => n10339, B => n1824, S => n1511, Z => n8298);
   U5498 : MUX2_X1 port map( A => n10340, B => n1813, S => n1511, Z => n8299);
   U5499 : MUX2_X1 port map( A => n10341, B => n1802, S => n1511, Z => n8300);
   U5500 : MUX2_X1 port map( A => n10278, B => n2949, S => n1512, Z => n8237);
   U5501 : MUX2_X1 port map( A => n10279, B => n2938, S => n1512, Z => n8238);
   U5502 : MUX2_X1 port map( A => n10280, B => n2927, S => n1512, Z => n8239);
   U5503 : MUX2_X1 port map( A => n10281, B => n2911, S => n1512, Z => n8240);
   U5504 : MUX2_X1 port map( A => n10282, B => n2900, S => n1512, Z => n8241);
   U5505 : MUX2_X1 port map( A => n10283, B => n2888, S => n1512, Z => n8242);
   U5506 : MUX2_X1 port map( A => n10284, B => n2877, S => n1512, Z => n8243);
   U5507 : MUX2_X1 port map( A => n10285, B => n2866, S => n1512, Z => n8244);
   U5508 : MUX2_X1 port map( A => n10286, B => n2855, S => n1512, Z => n8245);
   U5509 : MUX2_X1 port map( A => n10287, B => n2844, S => n1512, Z => n8246);
   U5510 : MUX2_X1 port map( A => n10288, B => n2833, S => n1512, Z => n8247);
   U5511 : MUX2_X1 port map( A => n10289, B => n2822, S => n1512, Z => n8248);
   U5512 : MUX2_X1 port map( A => n10290, B => n2811, S => n1513, Z => n8249);
   U5513 : MUX2_X1 port map( A => n10291, B => n2800, S => n1513, Z => n8250);
   U5514 : MUX2_X1 port map( A => n10292, B => n2789, S => n1513, Z => n8251);
   U5515 : MUX2_X1 port map( A => n10293, B => n2778, S => n1513, Z => n8252);
   U5516 : MUX2_X1 port map( A => n10294, B => n2767, S => n1513, Z => n8253);
   U5517 : MUX2_X1 port map( A => n10295, B => n2756, S => n1513, Z => n8254);
   U5518 : MUX2_X1 port map( A => n10296, B => n2745, S => n1513, Z => n8255);
   U5519 : MUX2_X1 port map( A => n10297, B => n2734, S => n1513, Z => n8256);
   U5520 : MUX2_X1 port map( A => n10298, B => n2723, S => n1513, Z => n8257);
   U5521 : MUX2_X1 port map( A => n10299, B => n2712, S => n1513, Z => n8258);
   U5522 : MUX2_X1 port map( A => n10300, B => n2605, S => n1513, Z => n8259);
   U5523 : MUX2_X1 port map( A => n10301, B => n2594, S => n1513, Z => n8260);
   U5524 : MUX2_X1 port map( A => n10302, B => n2583, S => n1514, Z => n8261);
   U5525 : MUX2_X1 port map( A => n10303, B => n2572, S => n1514, Z => n8262);
   U5526 : MUX2_X1 port map( A => n10304, B => n2561, S => n1514, Z => n8263);
   U5527 : MUX2_X1 port map( A => n10305, B => n2550, S => n1514, Z => n8264);
   U5528 : MUX2_X1 port map( A => n10306, B => n1835, S => n1514, Z => n8265);
   U5529 : MUX2_X1 port map( A => n10307, B => n1824, S => n1514, Z => n8266);
   U5530 : MUX2_X1 port map( A => n10308, B => n1813, S => n1514, Z => n8267);
   U5531 : MUX2_X1 port map( A => n10309, B => n1802, S => n1514, Z => n8268);
   U5532 : MUX2_X1 port map( A => n10246, B => n2949, S => n1515, Z => n8205);
   U5533 : MUX2_X1 port map( A => n10247, B => n2938, S => n1515, Z => n8206);
   U5534 : MUX2_X1 port map( A => n10248, B => n2927, S => n1515, Z => n8207);
   U5535 : MUX2_X1 port map( A => n10249, B => n2911, S => n1515, Z => n8208);
   U5536 : MUX2_X1 port map( A => n10250, B => n2900, S => n1515, Z => n8209);
   U5537 : MUX2_X1 port map( A => n10251, B => n2888, S => n1515, Z => n8210);
   U5538 : MUX2_X1 port map( A => n10252, B => n2877, S => n1515, Z => n8211);
   U5539 : MUX2_X1 port map( A => n10253, B => n2866, S => n1515, Z => n8212);
   U5540 : MUX2_X1 port map( A => n10254, B => n2855, S => n1515, Z => n8213);
   U5541 : MUX2_X1 port map( A => n10255, B => n2844, S => n1515, Z => n8214);
   U5542 : MUX2_X1 port map( A => n10256, B => n2833, S => n1515, Z => n8215);
   U5543 : MUX2_X1 port map( A => n10257, B => n2822, S => n1515, Z => n8216);
   U5544 : MUX2_X1 port map( A => n10258, B => n2811, S => n1516, Z => n8217);
   U5545 : MUX2_X1 port map( A => n10259, B => n2800, S => n1516, Z => n8218);
   U5546 : MUX2_X1 port map( A => n10260, B => n2789, S => n1516, Z => n8219);
   U5547 : MUX2_X1 port map( A => n10261, B => n2778, S => n1516, Z => n8220);
   U5548 : MUX2_X1 port map( A => n10262, B => n2767, S => n1516, Z => n8221);
   U5549 : MUX2_X1 port map( A => n10263, B => n2756, S => n1516, Z => n8222);
   U5550 : MUX2_X1 port map( A => n10264, B => n2745, S => n1516, Z => n8223);
   U5551 : MUX2_X1 port map( A => n10265, B => n2734, S => n1516, Z => n8224);
   U5552 : MUX2_X1 port map( A => n10266, B => n2723, S => n1516, Z => n8225);
   U5553 : MUX2_X1 port map( A => n10267, B => n2712, S => n1516, Z => n8226);
   U5554 : MUX2_X1 port map( A => n10268, B => n2605, S => n1516, Z => n8227);
   U5555 : MUX2_X1 port map( A => n10269, B => n2594, S => n1516, Z => n8228);
   U5556 : MUX2_X1 port map( A => n10270, B => n2583, S => n1517, Z => n8229);
   U5557 : MUX2_X1 port map( A => n10271, B => n2572, S => n1517, Z => n8230);
   U5558 : MUX2_X1 port map( A => n10272, B => n2561, S => n1517, Z => n8231);
   U5559 : MUX2_X1 port map( A => n10273, B => n2550, S => n1517, Z => n8232);
   U5560 : MUX2_X1 port map( A => n10274, B => n1835, S => n1517, Z => n8233);
   U5561 : MUX2_X1 port map( A => n10275, B => n1824, S => n1517, Z => n8234);
   U5562 : MUX2_X1 port map( A => n10276, B => n1813, S => n1517, Z => n8235);
   U5563 : MUX2_X1 port map( A => n10277, B => n1802, S => n1517, Z => n8236);
   U5564 : MUX2_X1 port map( A => n10214, B => n2949, S => n1518, Z => n8173);
   U5565 : MUX2_X1 port map( A => n10215, B => n2938, S => n1518, Z => n8174);
   U5566 : MUX2_X1 port map( A => n10216, B => n2927, S => n1518, Z => n8175);
   U5567 : MUX2_X1 port map( A => n10217, B => n2911, S => n1518, Z => n8176);
   U5568 : MUX2_X1 port map( A => n10218, B => n2900, S => n1518, Z => n8177);
   U5569 : MUX2_X1 port map( A => n10219, B => n2888, S => n1518, Z => n8178);
   U5570 : MUX2_X1 port map( A => n10220, B => n2877, S => n1518, Z => n8179);
   U5571 : MUX2_X1 port map( A => n10221, B => n2866, S => n1518, Z => n8180);
   U5572 : MUX2_X1 port map( A => n10222, B => n2855, S => n1518, Z => n8181);
   U5573 : MUX2_X1 port map( A => n10223, B => n2844, S => n1518, Z => n8182);
   U5574 : MUX2_X1 port map( A => n10224, B => n2833, S => n1518, Z => n8183);
   U5575 : MUX2_X1 port map( A => n10225, B => n2822, S => n1518, Z => n8184);
   U5576 : MUX2_X1 port map( A => n10226, B => n2811, S => n1519, Z => n8185);
   U5577 : MUX2_X1 port map( A => n10227, B => n2800, S => n1519, Z => n8186);
   U5578 : MUX2_X1 port map( A => n10228, B => n2789, S => n1519, Z => n8187);
   U5579 : MUX2_X1 port map( A => n10229, B => n2778, S => n1519, Z => n8188);
   U5580 : MUX2_X1 port map( A => n10230, B => n2767, S => n1519, Z => n8189);
   U5581 : MUX2_X1 port map( A => n10231, B => n2756, S => n1519, Z => n8190);
   U5582 : MUX2_X1 port map( A => n10232, B => n2745, S => n1519, Z => n8191);
   U5583 : MUX2_X1 port map( A => n10233, B => n2734, S => n1519, Z => n8192);
   U5584 : MUX2_X1 port map( A => n10234, B => n2723, S => n1519, Z => n8193);
   U5585 : MUX2_X1 port map( A => n10235, B => n2712, S => n1519, Z => n8194);
   U5586 : MUX2_X1 port map( A => n10236, B => n2605, S => n1519, Z => n8195);
   U5587 : MUX2_X1 port map( A => n10237, B => n2594, S => n1519, Z => n8196);
   U5588 : MUX2_X1 port map( A => n10238, B => n2583, S => n1520, Z => n8197);
   U5589 : MUX2_X1 port map( A => n10239, B => n2572, S => n1520, Z => n8198);
   U5590 : MUX2_X1 port map( A => n10240, B => n2561, S => n1520, Z => n8199);
   U5591 : MUX2_X1 port map( A => n10241, B => n2550, S => n1520, Z => n8200);
   U5592 : MUX2_X1 port map( A => n10242, B => n1835, S => n1520, Z => n8201);
   U5593 : MUX2_X1 port map( A => n10243, B => n1824, S => n1520, Z => n8202);
   U5594 : MUX2_X1 port map( A => n10244, B => n1813, S => n1520, Z => n8203);
   U5595 : MUX2_X1 port map( A => n10245, B => n1802, S => n1520, Z => n8204);
   U5596 : MUX2_X1 port map( A => n10182, B => n2949, S => n1521, Z => n8141);
   U5597 : MUX2_X1 port map( A => n10183, B => n2938, S => n1521, Z => n8142);
   U5598 : MUX2_X1 port map( A => n10184, B => n2927, S => n1521, Z => n8143);
   U5599 : MUX2_X1 port map( A => n10185, B => n2911, S => n1521, Z => n8144);
   U5600 : MUX2_X1 port map( A => n10186, B => n2900, S => n1521, Z => n8145);
   U5601 : MUX2_X1 port map( A => n10187, B => n2888, S => n1521, Z => n8146);
   U5602 : MUX2_X1 port map( A => n10188, B => n2877, S => n1521, Z => n8147);
   U5603 : MUX2_X1 port map( A => n10189, B => n2866, S => n1521, Z => n8148);
   U5604 : MUX2_X1 port map( A => n10190, B => n2855, S => n1521, Z => n8149);
   U5605 : MUX2_X1 port map( A => n10191, B => n2844, S => n1521, Z => n8150);
   U5606 : MUX2_X1 port map( A => n10192, B => n2833, S => n1521, Z => n8151);
   U5607 : MUX2_X1 port map( A => n10193, B => n2822, S => n1521, Z => n8152);
   U5608 : MUX2_X1 port map( A => n10194, B => n2811, S => n1522, Z => n8153);
   U5609 : MUX2_X1 port map( A => n10195, B => n2800, S => n1522, Z => n8154);
   U5610 : MUX2_X1 port map( A => n10196, B => n2789, S => n1522, Z => n8155);
   U5611 : MUX2_X1 port map( A => n10197, B => n2778, S => n1522, Z => n8156);
   U5612 : MUX2_X1 port map( A => n10198, B => n2767, S => n1522, Z => n8157);
   U5613 : MUX2_X1 port map( A => n10199, B => n2756, S => n1522, Z => n8158);
   U5614 : MUX2_X1 port map( A => n10200, B => n2745, S => n1522, Z => n8159);
   U5615 : MUX2_X1 port map( A => n10201, B => n2734, S => n1522, Z => n8160);
   U5616 : MUX2_X1 port map( A => n10202, B => n2723, S => n1522, Z => n8161);
   U5617 : MUX2_X1 port map( A => n10203, B => n2712, S => n1522, Z => n8162);
   U5618 : MUX2_X1 port map( A => n10204, B => n2605, S => n1522, Z => n8163);
   U5619 : MUX2_X1 port map( A => n10205, B => n2594, S => n1522, Z => n8164);
   U5620 : MUX2_X1 port map( A => n10206, B => n2583, S => n1523, Z => n8165);
   U5621 : MUX2_X1 port map( A => n10207, B => n2572, S => n1523, Z => n8166);
   U5622 : MUX2_X1 port map( A => n10208, B => n2561, S => n1523, Z => n8167);
   U5623 : MUX2_X1 port map( A => n10209, B => n2550, S => n1523, Z => n8168);
   U5624 : MUX2_X1 port map( A => n10210, B => n1835, S => n1523, Z => n8169);
   U5625 : MUX2_X1 port map( A => n10211, B => n1824, S => n1523, Z => n8170);
   U5626 : MUX2_X1 port map( A => n10212, B => n1813, S => n1523, Z => n8171);
   U5627 : MUX2_X1 port map( A => n10213, B => n1802, S => n1523, Z => n8172);
   U5628 : MUX2_X1 port map( A => n10150, B => n2949, S => n1524, Z => n8109);
   U5629 : MUX2_X1 port map( A => n10151, B => n2938, S => n1524, Z => n8110);
   U5630 : MUX2_X1 port map( A => n10152, B => n2927, S => n1524, Z => n8111);
   U5631 : MUX2_X1 port map( A => n10153, B => n2911, S => n1524, Z => n8112);
   U5632 : MUX2_X1 port map( A => n10154, B => n2900, S => n1524, Z => n8113);
   U5633 : MUX2_X1 port map( A => n10155, B => n2888, S => n1524, Z => n8114);
   U5634 : MUX2_X1 port map( A => n10156, B => n2877, S => n1524, Z => n8115);
   U5635 : MUX2_X1 port map( A => n10157, B => n2866, S => n1524, Z => n8116);
   U5636 : MUX2_X1 port map( A => n10158, B => n2855, S => n1524, Z => n8117);
   U5637 : MUX2_X1 port map( A => n10159, B => n2844, S => n1524, Z => n8118);
   U5638 : MUX2_X1 port map( A => n10160, B => n2833, S => n1524, Z => n8119);
   U5639 : MUX2_X1 port map( A => n10161, B => n2822, S => n1524, Z => n8120);
   U5640 : MUX2_X1 port map( A => n10162, B => n2811, S => n1525, Z => n8121);
   U5641 : MUX2_X1 port map( A => n10163, B => n2800, S => n1525, Z => n8122);
   U5642 : MUX2_X1 port map( A => n10164, B => n2789, S => n1525, Z => n8123);
   U5643 : MUX2_X1 port map( A => n10165, B => n2778, S => n1525, Z => n8124);
   U5644 : MUX2_X1 port map( A => n10166, B => n2767, S => n1525, Z => n8125);
   U5645 : MUX2_X1 port map( A => n10167, B => n2756, S => n1525, Z => n8126);
   U5646 : MUX2_X1 port map( A => n10168, B => n2745, S => n1525, Z => n8127);
   U5647 : MUX2_X1 port map( A => n10169, B => n2734, S => n1525, Z => n8128);
   U5648 : MUX2_X1 port map( A => n10170, B => n2723, S => n1525, Z => n8129);
   U5649 : MUX2_X1 port map( A => n10171, B => n2712, S => n1525, Z => n8130);
   U5650 : MUX2_X1 port map( A => n10172, B => n2605, S => n1525, Z => n8131);
   U5651 : MUX2_X1 port map( A => n10173, B => n2594, S => n1525, Z => n8132);
   U5652 : MUX2_X1 port map( A => n10174, B => n2583, S => n1526, Z => n8133);
   U5653 : MUX2_X1 port map( A => n10175, B => n2572, S => n1526, Z => n8134);
   U5654 : MUX2_X1 port map( A => n10176, B => n2561, S => n1526, Z => n8135);
   U5655 : MUX2_X1 port map( A => n10177, B => n2550, S => n1526, Z => n8136);
   U5656 : MUX2_X1 port map( A => n10178, B => n1835, S => n1526, Z => n8137);
   U5657 : MUX2_X1 port map( A => n10179, B => n1824, S => n1526, Z => n8138);
   U5658 : MUX2_X1 port map( A => n10180, B => n1813, S => n1526, Z => n8139);
   U5659 : MUX2_X1 port map( A => n10181, B => n1802, S => n1526, Z => n8140);
   U5660 : MUX2_X1 port map( A => n10118, B => n2949, S => n1527, Z => n8077);
   U5661 : MUX2_X1 port map( A => n10119, B => n2938, S => n1527, Z => n8078);
   U5662 : MUX2_X1 port map( A => n10120, B => n2927, S => n1527, Z => n8079);
   U5663 : MUX2_X1 port map( A => n10121, B => n2911, S => n1527, Z => n8080);
   U5664 : MUX2_X1 port map( A => n10122, B => n2900, S => n1527, Z => n8081);
   U5665 : MUX2_X1 port map( A => n10123, B => n2888, S => n1527, Z => n8082);
   U5666 : MUX2_X1 port map( A => n10124, B => n2877, S => n1527, Z => n8083);
   U5667 : MUX2_X1 port map( A => n10125, B => n2866, S => n1527, Z => n8084);
   U5668 : MUX2_X1 port map( A => n10126, B => n2855, S => n1527, Z => n8085);
   U5669 : MUX2_X1 port map( A => n10127, B => n2844, S => n1527, Z => n8086);
   U5670 : MUX2_X1 port map( A => n10128, B => n2833, S => n1527, Z => n8087);
   U5671 : MUX2_X1 port map( A => n10129, B => n2822, S => n1527, Z => n8088);
   U5672 : MUX2_X1 port map( A => n10130, B => n2811, S => n1528, Z => n8089);
   U5673 : MUX2_X1 port map( A => n10131, B => n2800, S => n1528, Z => n8090);
   U5674 : MUX2_X1 port map( A => n10132, B => n2789, S => n1528, Z => n8091);
   U5675 : MUX2_X1 port map( A => n10133, B => n2778, S => n1528, Z => n8092);
   U5676 : MUX2_X1 port map( A => n10134, B => n2767, S => n1528, Z => n8093);
   U5677 : MUX2_X1 port map( A => n10135, B => n2756, S => n1528, Z => n8094);
   U5678 : MUX2_X1 port map( A => n10136, B => n2745, S => n1528, Z => n8095);
   U5679 : MUX2_X1 port map( A => n10137, B => n2734, S => n1528, Z => n8096);
   U5680 : MUX2_X1 port map( A => n10138, B => n2723, S => n1528, Z => n8097);
   U5681 : MUX2_X1 port map( A => n10139, B => n2712, S => n1528, Z => n8098);
   U5682 : MUX2_X1 port map( A => n10140, B => n2605, S => n1528, Z => n8099);
   U5683 : MUX2_X1 port map( A => n10141, B => n2594, S => n1528, Z => n8100);
   U5684 : MUX2_X1 port map( A => n10142, B => n2583, S => n1529, Z => n8101);
   U5685 : MUX2_X1 port map( A => n10143, B => n2572, S => n1529, Z => n8102);
   U5686 : MUX2_X1 port map( A => n10144, B => n2561, S => n1529, Z => n8103);
   U5687 : MUX2_X1 port map( A => n10145, B => n2550, S => n1529, Z => n8104);
   U5688 : MUX2_X1 port map( A => n10146, B => n1835, S => n1529, Z => n8105);
   U5689 : MUX2_X1 port map( A => n10147, B => n1824, S => n1529, Z => n8106);
   U5690 : MUX2_X1 port map( A => n10148, B => n1813, S => n1529, Z => n8107);
   U5691 : MUX2_X1 port map( A => n10149, B => n1802, S => n1529, Z => n8108);
   U5692 : MUX2_X1 port map( A => REGISTERS_54_31_port, B => n2950, S => n1530,
                           Z => n8045);
   U5693 : MUX2_X1 port map( A => REGISTERS_54_30_port, B => n2939, S => n1530,
                           Z => n8046);
   U5694 : MUX2_X1 port map( A => REGISTERS_54_29_port, B => n2928, S => n1530,
                           Z => n8047);
   U5695 : MUX2_X1 port map( A => REGISTERS_54_28_port, B => n2912, S => n1530,
                           Z => n8048);
   U5696 : MUX2_X1 port map( A => REGISTERS_54_27_port, B => n2901, S => n1530,
                           Z => n8049);
   U5697 : MUX2_X1 port map( A => REGISTERS_54_26_port, B => n2889, S => n1530,
                           Z => n8050);
   U5698 : MUX2_X1 port map( A => REGISTERS_54_25_port, B => n2878, S => n1530,
                           Z => n8051);
   U5699 : MUX2_X1 port map( A => REGISTERS_54_24_port, B => n2867, S => n1530,
                           Z => n8052);
   U5700 : MUX2_X1 port map( A => REGISTERS_54_23_port, B => n2856, S => n1530,
                           Z => n8053);
   U5701 : MUX2_X1 port map( A => REGISTERS_54_22_port, B => n2845, S => n1530,
                           Z => n8054);
   U5702 : MUX2_X1 port map( A => REGISTERS_54_21_port, B => n2834, S => n1530,
                           Z => n8055);
   U5703 : MUX2_X1 port map( A => REGISTERS_54_20_port, B => n2823, S => n1530,
                           Z => n8056);
   U5704 : MUX2_X1 port map( A => REGISTERS_54_19_port, B => n2812, S => n1531,
                           Z => n8057);
   U5705 : MUX2_X1 port map( A => REGISTERS_54_18_port, B => n2801, S => n1531,
                           Z => n8058);
   U5706 : MUX2_X1 port map( A => REGISTERS_54_17_port, B => n2790, S => n1531,
                           Z => n8059);
   U5707 : MUX2_X1 port map( A => REGISTERS_54_16_port, B => n2779, S => n1531,
                           Z => n8060);
   U5708 : MUX2_X1 port map( A => REGISTERS_54_15_port, B => n2768, S => n1531,
                           Z => n8061);
   U5709 : MUX2_X1 port map( A => REGISTERS_54_14_port, B => n2757, S => n1531,
                           Z => n8062);
   U5710 : MUX2_X1 port map( A => REGISTERS_54_13_port, B => n2746, S => n1531,
                           Z => n8063);
   U5711 : MUX2_X1 port map( A => REGISTERS_54_12_port, B => n2735, S => n1531,
                           Z => n8064);
   U5712 : MUX2_X1 port map( A => REGISTERS_54_11_port, B => n2724, S => n1531,
                           Z => n8065);
   U5713 : MUX2_X1 port map( A => REGISTERS_54_10_port, B => n2713, S => n1531,
                           Z => n8066);
   U5714 : MUX2_X1 port map( A => REGISTERS_54_9_port, B => n2606, S => n1531, 
                           Z => n8067);
   U5715 : MUX2_X1 port map( A => REGISTERS_54_8_port, B => n2595, S => n1531, 
                           Z => n8068);
   U5716 : MUX2_X1 port map( A => REGISTERS_54_7_port, B => n2584, S => n1532, 
                           Z => n8069);
   U5717 : MUX2_X1 port map( A => REGISTERS_54_6_port, B => n2573, S => n1532, 
                           Z => n8070);
   U5718 : MUX2_X1 port map( A => REGISTERS_54_5_port, B => n2562, S => n1532, 
                           Z => n8071);
   U5719 : MUX2_X1 port map( A => REGISTERS_54_4_port, B => n2551, S => n1532, 
                           Z => n8072);
   U5720 : MUX2_X1 port map( A => REGISTERS_54_3_port, B => n1836, S => n1532, 
                           Z => n8073);
   U5721 : MUX2_X1 port map( A => REGISTERS_54_2_port, B => n1825, S => n1532, 
                           Z => n8074);
   U5722 : MUX2_X1 port map( A => REGISTERS_54_1_port, B => n1814, S => n1532, 
                           Z => n8075);
   U5723 : MUX2_X1 port map( A => REGISTERS_54_0_port, B => n1803, S => n1532, 
                           Z => n8076);
   U5724 : MUX2_X1 port map( A => REGISTERS_53_31_port, B => n2950, S => n1533,
                           Z => n8013);
   U5725 : MUX2_X1 port map( A => REGISTERS_53_30_port, B => n2939, S => n1533,
                           Z => n8014);
   U5726 : MUX2_X1 port map( A => REGISTERS_53_29_port, B => n2928, S => n1533,
                           Z => n8015);
   U5727 : MUX2_X1 port map( A => REGISTERS_53_28_port, B => n2912, S => n1533,
                           Z => n8016);
   U5728 : MUX2_X1 port map( A => REGISTERS_53_27_port, B => n2901, S => n1533,
                           Z => n8017);
   U5729 : MUX2_X1 port map( A => REGISTERS_53_26_port, B => n2889, S => n1533,
                           Z => n8018);
   U5730 : MUX2_X1 port map( A => REGISTERS_53_25_port, B => n2878, S => n1533,
                           Z => n8019);
   U5731 : MUX2_X1 port map( A => REGISTERS_53_24_port, B => n2867, S => n1533,
                           Z => n8020);
   U5732 : MUX2_X1 port map( A => REGISTERS_53_23_port, B => n2856, S => n1533,
                           Z => n8021);
   U5733 : MUX2_X1 port map( A => REGISTERS_53_22_port, B => n2845, S => n1533,
                           Z => n8022);
   U5734 : MUX2_X1 port map( A => REGISTERS_53_21_port, B => n2834, S => n1533,
                           Z => n8023);
   U5735 : MUX2_X1 port map( A => REGISTERS_53_20_port, B => n2823, S => n1533,
                           Z => n8024);
   U5736 : MUX2_X1 port map( A => REGISTERS_53_19_port, B => n2812, S => n1534,
                           Z => n8025);
   U5737 : MUX2_X1 port map( A => REGISTERS_53_18_port, B => n2801, S => n1534,
                           Z => n8026);
   U5738 : MUX2_X1 port map( A => REGISTERS_53_17_port, B => n2790, S => n1534,
                           Z => n8027);
   U5739 : MUX2_X1 port map( A => REGISTERS_53_16_port, B => n2779, S => n1534,
                           Z => n8028);
   U5740 : MUX2_X1 port map( A => REGISTERS_53_15_port, B => n2768, S => n1534,
                           Z => n8029);
   U5741 : MUX2_X1 port map( A => REGISTERS_53_14_port, B => n2757, S => n1534,
                           Z => n8030);
   U5742 : MUX2_X1 port map( A => REGISTERS_53_13_port, B => n2746, S => n1534,
                           Z => n8031);
   U5743 : MUX2_X1 port map( A => REGISTERS_53_12_port, B => n2735, S => n1534,
                           Z => n8032);
   U5744 : MUX2_X1 port map( A => REGISTERS_53_11_port, B => n2724, S => n1534,
                           Z => n8033);
   U5745 : MUX2_X1 port map( A => REGISTERS_53_10_port, B => n2713, S => n1534,
                           Z => n8034);
   U5746 : MUX2_X1 port map( A => REGISTERS_53_9_port, B => n2606, S => n1534, 
                           Z => n8035);
   U5747 : MUX2_X1 port map( A => REGISTERS_53_8_port, B => n2595, S => n1534, 
                           Z => n8036);
   U5748 : MUX2_X1 port map( A => REGISTERS_53_7_port, B => n2584, S => n1535, 
                           Z => n8037);
   U5749 : MUX2_X1 port map( A => REGISTERS_53_6_port, B => n2573, S => n1535, 
                           Z => n8038);
   U5750 : MUX2_X1 port map( A => REGISTERS_53_5_port, B => n2562, S => n1535, 
                           Z => n8039);
   U5751 : MUX2_X1 port map( A => REGISTERS_53_4_port, B => n2551, S => n1535, 
                           Z => n8040);
   U5752 : MUX2_X1 port map( A => REGISTERS_53_3_port, B => n1836, S => n1535, 
                           Z => n8041);
   U5753 : MUX2_X1 port map( A => REGISTERS_53_2_port, B => n1825, S => n1535, 
                           Z => n8042);
   U5754 : MUX2_X1 port map( A => REGISTERS_53_1_port, B => n1814, S => n1535, 
                           Z => n8043);
   U5755 : MUX2_X1 port map( A => REGISTERS_53_0_port, B => n1803, S => n1535, 
                           Z => n8044);
   U5756 : MUX2_X1 port map( A => REGISTERS_52_31_port, B => n2950, S => n1536,
                           Z => n7981);
   U5757 : MUX2_X1 port map( A => REGISTERS_52_30_port, B => n2939, S => n1536,
                           Z => n7982);
   U5758 : MUX2_X1 port map( A => REGISTERS_52_29_port, B => n2928, S => n1536,
                           Z => n7983);
   U5759 : MUX2_X1 port map( A => REGISTERS_52_28_port, B => n2912, S => n1536,
                           Z => n7984);
   U5760 : MUX2_X1 port map( A => REGISTERS_52_27_port, B => n2901, S => n1536,
                           Z => n7985);
   U5761 : MUX2_X1 port map( A => REGISTERS_52_26_port, B => n2889, S => n1536,
                           Z => n7986);
   U5762 : MUX2_X1 port map( A => REGISTERS_52_25_port, B => n2878, S => n1536,
                           Z => n7987);
   U5763 : MUX2_X1 port map( A => REGISTERS_52_24_port, B => n2867, S => n1536,
                           Z => n7988);
   U5764 : MUX2_X1 port map( A => REGISTERS_52_23_port, B => n2856, S => n1536,
                           Z => n7989);
   U5765 : MUX2_X1 port map( A => REGISTERS_52_22_port, B => n2845, S => n1536,
                           Z => n7990);
   U5766 : MUX2_X1 port map( A => REGISTERS_52_21_port, B => n2834, S => n1536,
                           Z => n7991);
   U5767 : MUX2_X1 port map( A => REGISTERS_52_20_port, B => n2823, S => n1536,
                           Z => n7992);
   U5768 : MUX2_X1 port map( A => REGISTERS_52_19_port, B => n2812, S => n1537,
                           Z => n7993);
   U5769 : MUX2_X1 port map( A => REGISTERS_52_18_port, B => n2801, S => n1537,
                           Z => n7994);
   U5770 : MUX2_X1 port map( A => REGISTERS_52_17_port, B => n2790, S => n1537,
                           Z => n7995);
   U5771 : MUX2_X1 port map( A => REGISTERS_52_16_port, B => n2779, S => n1537,
                           Z => n7996);
   U5772 : MUX2_X1 port map( A => REGISTERS_52_15_port, B => n2768, S => n1537,
                           Z => n7997);
   U5773 : MUX2_X1 port map( A => REGISTERS_52_14_port, B => n2757, S => n1537,
                           Z => n7998);
   U5774 : MUX2_X1 port map( A => REGISTERS_52_13_port, B => n2746, S => n1537,
                           Z => n7999);
   U5775 : MUX2_X1 port map( A => REGISTERS_52_12_port, B => n2735, S => n1537,
                           Z => n8000);
   U5776 : MUX2_X1 port map( A => REGISTERS_52_11_port, B => n2724, S => n1537,
                           Z => n8001);
   U5777 : MUX2_X1 port map( A => REGISTERS_52_10_port, B => n2713, S => n1537,
                           Z => n8002);
   U5778 : MUX2_X1 port map( A => REGISTERS_52_9_port, B => n2606, S => n1537, 
                           Z => n8003);
   U5779 : MUX2_X1 port map( A => REGISTERS_52_8_port, B => n2595, S => n1537, 
                           Z => n8004);
   U5780 : MUX2_X1 port map( A => REGISTERS_52_7_port, B => n2584, S => n1538, 
                           Z => n8005);
   U5781 : MUX2_X1 port map( A => REGISTERS_52_6_port, B => n2573, S => n1538, 
                           Z => n8006);
   U5782 : MUX2_X1 port map( A => REGISTERS_52_5_port, B => n2562, S => n1538, 
                           Z => n8007);
   U5783 : MUX2_X1 port map( A => REGISTERS_52_4_port, B => n2551, S => n1538, 
                           Z => n8008);
   U5784 : MUX2_X1 port map( A => REGISTERS_52_3_port, B => n1836, S => n1538, 
                           Z => n8009);
   U5785 : MUX2_X1 port map( A => REGISTERS_52_2_port, B => n1825, S => n1538, 
                           Z => n8010);
   U5786 : MUX2_X1 port map( A => REGISTERS_52_1_port, B => n1814, S => n1538, 
                           Z => n8011);
   U5787 : MUX2_X1 port map( A => REGISTERS_52_0_port, B => n1803, S => n1538, 
                           Z => n8012);
   U5788 : MUX2_X1 port map( A => REGISTERS_51_31_port, B => n2950, S => n1539,
                           Z => n7949);
   U5789 : MUX2_X1 port map( A => REGISTERS_51_30_port, B => n2939, S => n1539,
                           Z => n7950);
   U5790 : MUX2_X1 port map( A => REGISTERS_51_29_port, B => n2928, S => n1539,
                           Z => n7951);
   U5791 : MUX2_X1 port map( A => REGISTERS_51_28_port, B => n2912, S => n1539,
                           Z => n7952);
   U5792 : MUX2_X1 port map( A => REGISTERS_51_27_port, B => n2901, S => n1539,
                           Z => n7953);
   U5793 : MUX2_X1 port map( A => REGISTERS_51_26_port, B => n2889, S => n1539,
                           Z => n7954);
   U5794 : MUX2_X1 port map( A => REGISTERS_51_25_port, B => n2878, S => n1539,
                           Z => n7955);
   U5795 : MUX2_X1 port map( A => REGISTERS_51_24_port, B => n2867, S => n1539,
                           Z => n7956);
   U5796 : MUX2_X1 port map( A => REGISTERS_51_23_port, B => n2856, S => n1539,
                           Z => n7957);
   U5797 : MUX2_X1 port map( A => REGISTERS_51_22_port, B => n2845, S => n1539,
                           Z => n7958);
   U5798 : MUX2_X1 port map( A => REGISTERS_51_21_port, B => n2834, S => n1539,
                           Z => n7959);
   U5799 : MUX2_X1 port map( A => REGISTERS_51_20_port, B => n2823, S => n1539,
                           Z => n7960);
   U5800 : MUX2_X1 port map( A => REGISTERS_51_19_port, B => n2812, S => n1540,
                           Z => n7961);
   U5801 : MUX2_X1 port map( A => REGISTERS_51_18_port, B => n2801, S => n1540,
                           Z => n7962);
   U5802 : MUX2_X1 port map( A => REGISTERS_51_17_port, B => n2790, S => n1540,
                           Z => n7963);
   U5803 : MUX2_X1 port map( A => REGISTERS_51_16_port, B => n2779, S => n1540,
                           Z => n7964);
   U5804 : MUX2_X1 port map( A => REGISTERS_51_15_port, B => n2768, S => n1540,
                           Z => n7965);
   U5805 : MUX2_X1 port map( A => REGISTERS_51_14_port, B => n2757, S => n1540,
                           Z => n7966);
   U5806 : MUX2_X1 port map( A => REGISTERS_51_13_port, B => n2746, S => n1540,
                           Z => n7967);
   U5807 : MUX2_X1 port map( A => REGISTERS_51_12_port, B => n2735, S => n1540,
                           Z => n7968);
   U5808 : MUX2_X1 port map( A => REGISTERS_51_11_port, B => n2724, S => n1540,
                           Z => n7969);
   U5809 : MUX2_X1 port map( A => REGISTERS_51_10_port, B => n2713, S => n1540,
                           Z => n7970);
   U5810 : MUX2_X1 port map( A => REGISTERS_51_9_port, B => n2606, S => n1540, 
                           Z => n7971);
   U5811 : MUX2_X1 port map( A => REGISTERS_51_8_port, B => n2595, S => n1540, 
                           Z => n7972);
   U5812 : MUX2_X1 port map( A => REGISTERS_51_7_port, B => n2584, S => n1541, 
                           Z => n7973);
   U5813 : MUX2_X1 port map( A => REGISTERS_51_6_port, B => n2573, S => n1541, 
                           Z => n7974);
   U5814 : MUX2_X1 port map( A => REGISTERS_51_5_port, B => n2562, S => n1541, 
                           Z => n7975);
   U5815 : MUX2_X1 port map( A => REGISTERS_51_4_port, B => n2551, S => n1541, 
                           Z => n7976);
   U5816 : MUX2_X1 port map( A => REGISTERS_51_3_port, B => n1836, S => n1541, 
                           Z => n7977);
   U5817 : MUX2_X1 port map( A => REGISTERS_51_2_port, B => n1825, S => n1541, 
                           Z => n7978);
   U5818 : MUX2_X1 port map( A => REGISTERS_51_1_port, B => n1814, S => n1541, 
                           Z => n7979);
   U5819 : MUX2_X1 port map( A => REGISTERS_51_0_port, B => n1803, S => n1541, 
                           Z => n7980);
   U5820 : MUX2_X1 port map( A => REGISTERS_50_31_port, B => n2950, S => n1542,
                           Z => n7917);
   U5821 : MUX2_X1 port map( A => REGISTERS_50_30_port, B => n2939, S => n1542,
                           Z => n7918);
   U5822 : MUX2_X1 port map( A => REGISTERS_50_29_port, B => n2928, S => n1542,
                           Z => n7919);
   U5823 : MUX2_X1 port map( A => REGISTERS_50_28_port, B => n2912, S => n1542,
                           Z => n7920);
   U5824 : MUX2_X1 port map( A => REGISTERS_50_27_port, B => n2901, S => n1542,
                           Z => n7921);
   U5825 : MUX2_X1 port map( A => REGISTERS_50_26_port, B => n2889, S => n1542,
                           Z => n7922);
   U5826 : MUX2_X1 port map( A => REGISTERS_50_25_port, B => n2878, S => n1542,
                           Z => n7923);
   U5827 : MUX2_X1 port map( A => REGISTERS_50_24_port, B => n2867, S => n1542,
                           Z => n7924);
   U5828 : MUX2_X1 port map( A => REGISTERS_50_23_port, B => n2856, S => n1542,
                           Z => n7925);
   U5829 : MUX2_X1 port map( A => REGISTERS_50_22_port, B => n2845, S => n1542,
                           Z => n7926);
   U5830 : MUX2_X1 port map( A => REGISTERS_50_21_port, B => n2834, S => n1542,
                           Z => n7927);
   U5831 : MUX2_X1 port map( A => REGISTERS_50_20_port, B => n2823, S => n1542,
                           Z => n7928);
   U5832 : MUX2_X1 port map( A => REGISTERS_50_19_port, B => n2812, S => n1543,
                           Z => n7929);
   U5833 : MUX2_X1 port map( A => REGISTERS_50_18_port, B => n2801, S => n1543,
                           Z => n7930);
   U5834 : MUX2_X1 port map( A => REGISTERS_50_17_port, B => n2790, S => n1543,
                           Z => n7931);
   U5835 : MUX2_X1 port map( A => REGISTERS_50_16_port, B => n2779, S => n1543,
                           Z => n7932);
   U5836 : MUX2_X1 port map( A => REGISTERS_50_15_port, B => n2768, S => n1543,
                           Z => n7933);
   U5837 : MUX2_X1 port map( A => REGISTERS_50_14_port, B => n2757, S => n1543,
                           Z => n7934);
   U5838 : MUX2_X1 port map( A => REGISTERS_50_13_port, B => n2746, S => n1543,
                           Z => n7935);
   U5839 : MUX2_X1 port map( A => REGISTERS_50_12_port, B => n2735, S => n1543,
                           Z => n7936);
   U5840 : MUX2_X1 port map( A => REGISTERS_50_11_port, B => n2724, S => n1543,
                           Z => n7937);
   U5841 : MUX2_X1 port map( A => REGISTERS_50_10_port, B => n2713, S => n1543,
                           Z => n7938);
   U5842 : MUX2_X1 port map( A => REGISTERS_50_9_port, B => n2606, S => n1543, 
                           Z => n7939);
   U5843 : MUX2_X1 port map( A => REGISTERS_50_8_port, B => n2595, S => n1543, 
                           Z => n7940);
   U5844 : MUX2_X1 port map( A => REGISTERS_50_7_port, B => n2584, S => n1544, 
                           Z => n7941);
   U5845 : MUX2_X1 port map( A => REGISTERS_50_6_port, B => n2573, S => n1544, 
                           Z => n7942);
   U5846 : MUX2_X1 port map( A => REGISTERS_50_5_port, B => n2562, S => n1544, 
                           Z => n7943);
   U5847 : MUX2_X1 port map( A => REGISTERS_50_4_port, B => n2551, S => n1544, 
                           Z => n7944);
   U5848 : MUX2_X1 port map( A => REGISTERS_50_3_port, B => n1836, S => n1544, 
                           Z => n7945);
   U5849 : MUX2_X1 port map( A => REGISTERS_50_2_port, B => n1825, S => n1544, 
                           Z => n7946);
   U5850 : MUX2_X1 port map( A => REGISTERS_50_1_port, B => n1814, S => n1544, 
                           Z => n7947);
   U5851 : MUX2_X1 port map( A => REGISTERS_50_0_port, B => n1803, S => n1544, 
                           Z => n7948);
   U5852 : MUX2_X1 port map( A => REGISTERS_49_31_port, B => n2950, S => n1545,
                           Z => n7885);
   U5853 : MUX2_X1 port map( A => REGISTERS_49_30_port, B => n2939, S => n1545,
                           Z => n7886);
   U5854 : MUX2_X1 port map( A => REGISTERS_49_29_port, B => n2928, S => n1545,
                           Z => n7887);
   U5855 : MUX2_X1 port map( A => REGISTERS_49_28_port, B => n2912, S => n1545,
                           Z => n7888);
   U5856 : MUX2_X1 port map( A => REGISTERS_49_27_port, B => n2901, S => n1545,
                           Z => n7889);
   U5857 : MUX2_X1 port map( A => REGISTERS_49_26_port, B => n2889, S => n1545,
                           Z => n7890);
   U5858 : MUX2_X1 port map( A => REGISTERS_49_25_port, B => n2878, S => n1545,
                           Z => n7891);
   U5859 : MUX2_X1 port map( A => REGISTERS_49_24_port, B => n2867, S => n1545,
                           Z => n7892);
   U5860 : MUX2_X1 port map( A => REGISTERS_49_23_port, B => n2856, S => n1545,
                           Z => n7893);
   U5861 : MUX2_X1 port map( A => REGISTERS_49_22_port, B => n2845, S => n1545,
                           Z => n7894);
   U5862 : MUX2_X1 port map( A => REGISTERS_49_21_port, B => n2834, S => n1545,
                           Z => n7895);
   U5863 : MUX2_X1 port map( A => REGISTERS_49_20_port, B => n2823, S => n1545,
                           Z => n7896);
   U5864 : MUX2_X1 port map( A => REGISTERS_49_19_port, B => n2812, S => n1546,
                           Z => n7897);
   U5865 : MUX2_X1 port map( A => REGISTERS_49_18_port, B => n2801, S => n1546,
                           Z => n7898);
   U5866 : MUX2_X1 port map( A => REGISTERS_49_17_port, B => n2790, S => n1546,
                           Z => n7899);
   U5867 : MUX2_X1 port map( A => REGISTERS_49_16_port, B => n2779, S => n1546,
                           Z => n7900);
   U5868 : MUX2_X1 port map( A => REGISTERS_49_15_port, B => n2768, S => n1546,
                           Z => n7901);
   U5869 : MUX2_X1 port map( A => REGISTERS_49_14_port, B => n2757, S => n1546,
                           Z => n7902);
   U5870 : MUX2_X1 port map( A => REGISTERS_49_13_port, B => n2746, S => n1546,
                           Z => n7903);
   U5871 : MUX2_X1 port map( A => REGISTERS_49_12_port, B => n2735, S => n1546,
                           Z => n7904);
   U5872 : MUX2_X1 port map( A => REGISTERS_49_11_port, B => n2724, S => n1546,
                           Z => n7905);
   U5873 : MUX2_X1 port map( A => REGISTERS_49_10_port, B => n2713, S => n1546,
                           Z => n7906);
   U5874 : MUX2_X1 port map( A => REGISTERS_49_9_port, B => n2606, S => n1546, 
                           Z => n7907);
   U5875 : MUX2_X1 port map( A => REGISTERS_49_8_port, B => n2595, S => n1546, 
                           Z => n7908);
   U5876 : MUX2_X1 port map( A => REGISTERS_49_7_port, B => n2584, S => n1547, 
                           Z => n7909);
   U5877 : MUX2_X1 port map( A => REGISTERS_49_6_port, B => n2573, S => n1547, 
                           Z => n7910);
   U5878 : MUX2_X1 port map( A => REGISTERS_49_5_port, B => n2562, S => n1547, 
                           Z => n7911);
   U5879 : MUX2_X1 port map( A => REGISTERS_49_4_port, B => n2551, S => n1547, 
                           Z => n7912);
   U5880 : MUX2_X1 port map( A => REGISTERS_49_3_port, B => n1836, S => n1547, 
                           Z => n7913);
   U5881 : MUX2_X1 port map( A => REGISTERS_49_2_port, B => n1825, S => n1547, 
                           Z => n7914);
   U5882 : MUX2_X1 port map( A => REGISTERS_49_1_port, B => n1814, S => n1547, 
                           Z => n7915);
   U5883 : MUX2_X1 port map( A => REGISTERS_49_0_port, B => n1803, S => n1547, 
                           Z => n7916);
   U5884 : MUX2_X1 port map( A => n10086, B => n2950, S => n1548, Z => n7853);
   U5885 : MUX2_X1 port map( A => n10087, B => n2939, S => n1548, Z => n7854);
   U5886 : MUX2_X1 port map( A => n10088, B => n2928, S => n1548, Z => n7855);
   U5887 : MUX2_X1 port map( A => n10089, B => n2912, S => n1548, Z => n7856);
   U5888 : MUX2_X1 port map( A => n10090, B => n2901, S => n1548, Z => n7857);
   U5889 : MUX2_X1 port map( A => n10091, B => n2889, S => n1548, Z => n7858);
   U5890 : MUX2_X1 port map( A => n10092, B => n2878, S => n1548, Z => n7859);
   U5891 : MUX2_X1 port map( A => n10093, B => n2867, S => n1548, Z => n7860);
   U5892 : MUX2_X1 port map( A => n10094, B => n2856, S => n1548, Z => n7861);
   U5893 : MUX2_X1 port map( A => n10095, B => n2845, S => n1548, Z => n7862);
   U5894 : MUX2_X1 port map( A => n10096, B => n2834, S => n1548, Z => n7863);
   U5895 : MUX2_X1 port map( A => n10097, B => n2823, S => n1548, Z => n7864);
   U5896 : MUX2_X1 port map( A => n10098, B => n2812, S => n1549, Z => n7865);
   U5897 : MUX2_X1 port map( A => n10099, B => n2801, S => n1549, Z => n7866);
   U5898 : MUX2_X1 port map( A => n10100, B => n2790, S => n1549, Z => n7867);
   U5899 : MUX2_X1 port map( A => n10101, B => n2779, S => n1549, Z => n7868);
   U5900 : MUX2_X1 port map( A => n10102, B => n2768, S => n1549, Z => n7869);
   U5901 : MUX2_X1 port map( A => n10103, B => n2757, S => n1549, Z => n7870);
   U5902 : MUX2_X1 port map( A => n10104, B => n2746, S => n1549, Z => n7871);
   U5903 : MUX2_X1 port map( A => n10105, B => n2735, S => n1549, Z => n7872);
   U5904 : MUX2_X1 port map( A => n10106, B => n2724, S => n1549, Z => n7873);
   U5905 : MUX2_X1 port map( A => n10107, B => n2713, S => n1549, Z => n7874);
   U5906 : MUX2_X1 port map( A => n10108, B => n2606, S => n1549, Z => n7875);
   U5907 : MUX2_X1 port map( A => n10109, B => n2595, S => n1549, Z => n7876);
   U5908 : MUX2_X1 port map( A => n10110, B => n2584, S => n1550, Z => n7877);
   U5909 : MUX2_X1 port map( A => n10111, B => n2573, S => n1550, Z => n7878);
   U5910 : MUX2_X1 port map( A => n10112, B => n2562, S => n1550, Z => n7879);
   U5911 : MUX2_X1 port map( A => n10113, B => n2551, S => n1550, Z => n7880);
   U5912 : MUX2_X1 port map( A => n10114, B => n1836, S => n1550, Z => n7881);
   U5913 : MUX2_X1 port map( A => n10115, B => n1825, S => n1550, Z => n7882);
   U5914 : MUX2_X1 port map( A => n10116, B => n1814, S => n1550, Z => n7883);
   U5915 : MUX2_X1 port map( A => n10117, B => n1803, S => n1550, Z => n7884);
   U5916 : MUX2_X1 port map( A => n10054, B => n2950, S => n1551, Z => n7821);
   U5917 : MUX2_X1 port map( A => n10055, B => n2939, S => n1551, Z => n7822);
   U5918 : MUX2_X1 port map( A => n10056, B => n2928, S => n1551, Z => n7823);
   U5919 : MUX2_X1 port map( A => n10057, B => n2912, S => n1551, Z => n7824);
   U5920 : MUX2_X1 port map( A => n10058, B => n2901, S => n1551, Z => n7825);
   U5921 : MUX2_X1 port map( A => n10059, B => n2889, S => n1551, Z => n7826);
   U5922 : MUX2_X1 port map( A => n10060, B => n2878, S => n1551, Z => n7827);
   U5923 : MUX2_X1 port map( A => n10061, B => n2867, S => n1551, Z => n7828);
   U5924 : MUX2_X1 port map( A => n10062, B => n2856, S => n1551, Z => n7829);
   U5925 : MUX2_X1 port map( A => n10063, B => n2845, S => n1551, Z => n7830);
   U5926 : MUX2_X1 port map( A => n10064, B => n2834, S => n1551, Z => n7831);
   U5927 : MUX2_X1 port map( A => n10065, B => n2823, S => n1551, Z => n7832);
   U5928 : MUX2_X1 port map( A => n10066, B => n2812, S => n1648, Z => n7833);
   U5929 : MUX2_X1 port map( A => n10067, B => n2801, S => n1648, Z => n7834);
   U5930 : MUX2_X1 port map( A => n10068, B => n2790, S => n1648, Z => n7835);
   U5931 : MUX2_X1 port map( A => n10069, B => n2779, S => n1648, Z => n7836);
   U5932 : MUX2_X1 port map( A => n10070, B => n2768, S => n1648, Z => n7837);
   U5933 : MUX2_X1 port map( A => n10071, B => n2757, S => n1648, Z => n7838);
   U5934 : MUX2_X1 port map( A => n10072, B => n2746, S => n1648, Z => n7839);
   U5935 : MUX2_X1 port map( A => n10073, B => n2735, S => n1648, Z => n7840);
   U5936 : MUX2_X1 port map( A => n10074, B => n2724, S => n1648, Z => n7841);
   U5937 : MUX2_X1 port map( A => n10075, B => n2713, S => n1648, Z => n7842);
   U5938 : MUX2_X1 port map( A => n10076, B => n2606, S => n1648, Z => n7843);
   U5939 : MUX2_X1 port map( A => n10077, B => n2595, S => n1648, Z => n7844);
   U5940 : MUX2_X1 port map( A => n10078, B => n2584, S => n1649, Z => n7845);
   U5941 : MUX2_X1 port map( A => n10079, B => n2573, S => n1649, Z => n7846);
   U5942 : MUX2_X1 port map( A => n10080, B => n2562, S => n1649, Z => n7847);
   U5943 : MUX2_X1 port map( A => n10081, B => n2551, S => n1649, Z => n7848);
   U5944 : MUX2_X1 port map( A => n10082, B => n1836, S => n1649, Z => n7849);
   U5945 : MUX2_X1 port map( A => n10083, B => n1825, S => n1649, Z => n7850);
   U5946 : MUX2_X1 port map( A => n10084, B => n1814, S => n1649, Z => n7851);
   U5947 : MUX2_X1 port map( A => n10085, B => n1803, S => n1649, Z => n7852);
   U5948 : MUX2_X1 port map( A => n10022, B => n2950, S => n1650, Z => n7789);
   U5949 : MUX2_X1 port map( A => n10023, B => n2939, S => n1650, Z => n7790);
   U5950 : MUX2_X1 port map( A => n10024, B => n2928, S => n1650, Z => n7791);
   U5951 : MUX2_X1 port map( A => n10025, B => n2912, S => n1650, Z => n7792);
   U5952 : MUX2_X1 port map( A => n10026, B => n2901, S => n1650, Z => n7793);
   U5953 : MUX2_X1 port map( A => n10027, B => n2889, S => n1650, Z => n7794);
   U5954 : MUX2_X1 port map( A => n10028, B => n2878, S => n1650, Z => n7795);
   U5955 : MUX2_X1 port map( A => n10029, B => n2867, S => n1650, Z => n7796);
   U5956 : MUX2_X1 port map( A => n10030, B => n2856, S => n1650, Z => n7797);
   U5957 : MUX2_X1 port map( A => n10031, B => n2845, S => n1650, Z => n7798);
   U5958 : MUX2_X1 port map( A => n10032, B => n2834, S => n1650, Z => n7799);
   U5959 : MUX2_X1 port map( A => n10033, B => n2823, S => n1650, Z => n7800);
   U5960 : MUX2_X1 port map( A => n10034, B => n2812, S => n1651, Z => n7801);
   U5961 : MUX2_X1 port map( A => n10035, B => n2801, S => n1651, Z => n7802);
   U5962 : MUX2_X1 port map( A => n10036, B => n2790, S => n1651, Z => n7803);
   U5963 : MUX2_X1 port map( A => n10037, B => n2779, S => n1651, Z => n7804);
   U5964 : MUX2_X1 port map( A => n10038, B => n2768, S => n1651, Z => n7805);
   U5965 : MUX2_X1 port map( A => n10039, B => n2757, S => n1651, Z => n7806);
   U5966 : MUX2_X1 port map( A => n10040, B => n2746, S => n1651, Z => n7807);
   U5967 : MUX2_X1 port map( A => n10041, B => n2735, S => n1651, Z => n7808);
   U5968 : MUX2_X1 port map( A => n10042, B => n2724, S => n1651, Z => n7809);
   U5969 : MUX2_X1 port map( A => n10043, B => n2713, S => n1651, Z => n7810);
   U5970 : MUX2_X1 port map( A => n10044, B => n2606, S => n1651, Z => n7811);
   U5971 : MUX2_X1 port map( A => n10045, B => n2595, S => n1651, Z => n7812);
   U5972 : MUX2_X1 port map( A => n10046, B => n2584, S => n1652, Z => n7813);
   U5973 : MUX2_X1 port map( A => n10047, B => n2573, S => n1652, Z => n7814);
   U5974 : MUX2_X1 port map( A => n10048, B => n2562, S => n1652, Z => n7815);
   U5975 : MUX2_X1 port map( A => n10049, B => n2551, S => n1652, Z => n7816);
   U5976 : MUX2_X1 port map( A => n10050, B => n1836, S => n1652, Z => n7817);
   U5977 : MUX2_X1 port map( A => n10051, B => n1825, S => n1652, Z => n7818);
   U5978 : MUX2_X1 port map( A => n10052, B => n1814, S => n1652, Z => n7819);
   U5979 : MUX2_X1 port map( A => n10053, B => n1803, S => n1652, Z => n7820);
   U5980 : MUX2_X1 port map( A => REGISTERS_45_31_port, B => n2950, S => n1653,
                           Z => n7757);
   U5981 : MUX2_X1 port map( A => REGISTERS_45_30_port, B => n2939, S => n1653,
                           Z => n7758);
   U5982 : MUX2_X1 port map( A => REGISTERS_45_29_port, B => n2928, S => n1653,
                           Z => n7759);
   U5983 : MUX2_X1 port map( A => REGISTERS_45_28_port, B => n2912, S => n1653,
                           Z => n7760);
   U5984 : MUX2_X1 port map( A => REGISTERS_45_27_port, B => n2901, S => n1653,
                           Z => n7761);
   U5985 : MUX2_X1 port map( A => REGISTERS_45_26_port, B => n2889, S => n1653,
                           Z => n7762);
   U5986 : MUX2_X1 port map( A => REGISTERS_45_25_port, B => n2878, S => n1653,
                           Z => n7763);
   U5987 : MUX2_X1 port map( A => REGISTERS_45_24_port, B => n2867, S => n1653,
                           Z => n7764);
   U5988 : MUX2_X1 port map( A => REGISTERS_45_23_port, B => n2856, S => n1653,
                           Z => n7765);
   U5989 : MUX2_X1 port map( A => REGISTERS_45_22_port, B => n2845, S => n1653,
                           Z => n7766);
   U5990 : MUX2_X1 port map( A => REGISTERS_45_21_port, B => n2834, S => n1653,
                           Z => n7767);
   U5991 : MUX2_X1 port map( A => REGISTERS_45_20_port, B => n2823, S => n1653,
                           Z => n7768);
   U5992 : MUX2_X1 port map( A => REGISTERS_45_19_port, B => n2812, S => n1654,
                           Z => n7769);
   U5993 : MUX2_X1 port map( A => REGISTERS_45_18_port, B => n2801, S => n1654,
                           Z => n7770);
   U5994 : MUX2_X1 port map( A => REGISTERS_45_17_port, B => n2790, S => n1654,
                           Z => n7771);
   U5995 : MUX2_X1 port map( A => REGISTERS_45_16_port, B => n2779, S => n1654,
                           Z => n7772);
   U5996 : MUX2_X1 port map( A => REGISTERS_45_15_port, B => n2768, S => n1654,
                           Z => n7773);
   U5997 : MUX2_X1 port map( A => REGISTERS_45_14_port, B => n2757, S => n1654,
                           Z => n7774);
   U5998 : MUX2_X1 port map( A => REGISTERS_45_13_port, B => n2746, S => n1654,
                           Z => n7775);
   U5999 : MUX2_X1 port map( A => REGISTERS_45_12_port, B => n2735, S => n1654,
                           Z => n7776);
   U6000 : MUX2_X1 port map( A => REGISTERS_45_11_port, B => n2724, S => n1654,
                           Z => n7777);
   U6001 : MUX2_X1 port map( A => REGISTERS_45_10_port, B => n2713, S => n1654,
                           Z => n7778);
   U6002 : MUX2_X1 port map( A => REGISTERS_45_9_port, B => n2606, S => n1654, 
                           Z => n7779);
   U6003 : MUX2_X1 port map( A => REGISTERS_45_8_port, B => n2595, S => n1654, 
                           Z => n7780);
   U6004 : MUX2_X1 port map( A => REGISTERS_45_7_port, B => n2584, S => n1655, 
                           Z => n7781);
   U6005 : MUX2_X1 port map( A => REGISTERS_45_6_port, B => n2573, S => n1655, 
                           Z => n7782);
   U6006 : MUX2_X1 port map( A => REGISTERS_45_5_port, B => n2562, S => n1655, 
                           Z => n7783);
   U6007 : MUX2_X1 port map( A => REGISTERS_45_4_port, B => n2551, S => n1655, 
                           Z => n7784);
   U6008 : MUX2_X1 port map( A => REGISTERS_45_3_port, B => n1836, S => n1655, 
                           Z => n7785);
   U6009 : MUX2_X1 port map( A => REGISTERS_45_2_port, B => n1825, S => n1655, 
                           Z => n7786);
   U6010 : MUX2_X1 port map( A => REGISTERS_45_1_port, B => n1814, S => n1655, 
                           Z => n7787);
   U6011 : MUX2_X1 port map( A => REGISTERS_45_0_port, B => n1803, S => n1655, 
                           Z => n7788);
   U6012 : MUX2_X1 port map( A => REGISTERS_44_31_port, B => n2950, S => n1656,
                           Z => n7725);
   U6013 : MUX2_X1 port map( A => REGISTERS_44_30_port, B => n2939, S => n1656,
                           Z => n7726);
   U6014 : MUX2_X1 port map( A => REGISTERS_44_29_port, B => n2928, S => n1656,
                           Z => n7727);
   U6015 : MUX2_X1 port map( A => REGISTERS_44_28_port, B => n2912, S => n1656,
                           Z => n7728);
   U6016 : MUX2_X1 port map( A => REGISTERS_44_27_port, B => n2901, S => n1656,
                           Z => n7729);
   U6017 : MUX2_X1 port map( A => REGISTERS_44_26_port, B => n2889, S => n1656,
                           Z => n7730);
   U6018 : MUX2_X1 port map( A => REGISTERS_44_25_port, B => n2878, S => n1656,
                           Z => n7731);
   U6019 : MUX2_X1 port map( A => REGISTERS_44_24_port, B => n2867, S => n1656,
                           Z => n7732);
   U6020 : MUX2_X1 port map( A => REGISTERS_44_23_port, B => n2856, S => n1656,
                           Z => n7733);
   U6021 : MUX2_X1 port map( A => REGISTERS_44_22_port, B => n2845, S => n1656,
                           Z => n7734);
   U6022 : MUX2_X1 port map( A => REGISTERS_44_21_port, B => n2834, S => n1656,
                           Z => n7735);
   U6023 : MUX2_X1 port map( A => REGISTERS_44_20_port, B => n2823, S => n1656,
                           Z => n7736);
   U6024 : MUX2_X1 port map( A => REGISTERS_44_19_port, B => n2812, S => n1657,
                           Z => n7737);
   U6025 : MUX2_X1 port map( A => REGISTERS_44_18_port, B => n2801, S => n1657,
                           Z => n7738);
   U6026 : MUX2_X1 port map( A => REGISTERS_44_17_port, B => n2790, S => n1657,
                           Z => n7739);
   U6027 : MUX2_X1 port map( A => REGISTERS_44_16_port, B => n2779, S => n1657,
                           Z => n7740);
   U6028 : MUX2_X1 port map( A => REGISTERS_44_15_port, B => n2768, S => n1657,
                           Z => n7741);
   U6029 : MUX2_X1 port map( A => REGISTERS_44_14_port, B => n2757, S => n1657,
                           Z => n7742);
   U6030 : MUX2_X1 port map( A => REGISTERS_44_13_port, B => n2746, S => n1657,
                           Z => n7743);
   U6031 : MUX2_X1 port map( A => REGISTERS_44_12_port, B => n2735, S => n1657,
                           Z => n7744);
   U6032 : MUX2_X1 port map( A => REGISTERS_44_11_port, B => n2724, S => n1657,
                           Z => n7745);
   U6033 : MUX2_X1 port map( A => REGISTERS_44_10_port, B => n2713, S => n1657,
                           Z => n7746);
   U6034 : MUX2_X1 port map( A => REGISTERS_44_9_port, B => n2606, S => n1657, 
                           Z => n7747);
   U6035 : MUX2_X1 port map( A => REGISTERS_44_8_port, B => n2595, S => n1657, 
                           Z => n7748);
   U6036 : MUX2_X1 port map( A => REGISTERS_44_7_port, B => n2584, S => n1658, 
                           Z => n7749);
   U6037 : MUX2_X1 port map( A => REGISTERS_44_6_port, B => n2573, S => n1658, 
                           Z => n7750);
   U6038 : MUX2_X1 port map( A => REGISTERS_44_5_port, B => n2562, S => n1658, 
                           Z => n7751);
   U6039 : MUX2_X1 port map( A => REGISTERS_44_4_port, B => n2551, S => n1658, 
                           Z => n7752);
   U6040 : MUX2_X1 port map( A => REGISTERS_44_3_port, B => n1836, S => n1658, 
                           Z => n7753);
   U6041 : MUX2_X1 port map( A => REGISTERS_44_2_port, B => n1825, S => n1658, 
                           Z => n7754);
   U6042 : MUX2_X1 port map( A => REGISTERS_44_1_port, B => n1814, S => n1658, 
                           Z => n7755);
   U6043 : MUX2_X1 port map( A => REGISTERS_44_0_port, B => n1803, S => n1658, 
                           Z => n7756);
   U6044 : MUX2_X1 port map( A => REGISTERS_43_31_port, B => n2951, S => n1659,
                           Z => n7693);
   U6045 : MUX2_X1 port map( A => REGISTERS_43_30_port, B => n2940, S => n1659,
                           Z => n7694);
   U6046 : MUX2_X1 port map( A => REGISTERS_43_29_port, B => n2929, S => n1659,
                           Z => n7695);
   U6047 : MUX2_X1 port map( A => REGISTERS_43_28_port, B => n2913, S => n1659,
                           Z => n7696);
   U6048 : MUX2_X1 port map( A => REGISTERS_43_27_port, B => n2902, S => n1659,
                           Z => n7697);
   U6049 : MUX2_X1 port map( A => REGISTERS_43_26_port, B => n2890, S => n1659,
                           Z => n7698);
   U6050 : MUX2_X1 port map( A => REGISTERS_43_25_port, B => n2879, S => n1659,
                           Z => n7699);
   U6051 : MUX2_X1 port map( A => REGISTERS_43_24_port, B => n2868, S => n1659,
                           Z => n7700);
   U6052 : MUX2_X1 port map( A => REGISTERS_43_23_port, B => n2857, S => n1659,
                           Z => n7701);
   U6053 : MUX2_X1 port map( A => REGISTERS_43_22_port, B => n2846, S => n1659,
                           Z => n7702);
   U6054 : MUX2_X1 port map( A => REGISTERS_43_21_port, B => n2835, S => n1659,
                           Z => n7703);
   U6055 : MUX2_X1 port map( A => REGISTERS_43_20_port, B => n2824, S => n1659,
                           Z => n7704);
   U6056 : MUX2_X1 port map( A => REGISTERS_43_19_port, B => n2813, S => n1660,
                           Z => n7705);
   U6057 : MUX2_X1 port map( A => REGISTERS_43_18_port, B => n2802, S => n1660,
                           Z => n7706);
   U6058 : MUX2_X1 port map( A => REGISTERS_43_17_port, B => n2791, S => n1660,
                           Z => n7707);
   U6059 : MUX2_X1 port map( A => REGISTERS_43_16_port, B => n2780, S => n1660,
                           Z => n7708);
   U6060 : MUX2_X1 port map( A => REGISTERS_43_15_port, B => n2769, S => n1660,
                           Z => n7709);
   U6061 : MUX2_X1 port map( A => REGISTERS_43_14_port, B => n2758, S => n1660,
                           Z => n7710);
   U6062 : MUX2_X1 port map( A => REGISTERS_43_13_port, B => n2747, S => n1660,
                           Z => n7711);
   U6063 : MUX2_X1 port map( A => REGISTERS_43_12_port, B => n2736, S => n1660,
                           Z => n7712);
   U6064 : MUX2_X1 port map( A => REGISTERS_43_11_port, B => n2725, S => n1660,
                           Z => n7713);
   U6065 : MUX2_X1 port map( A => REGISTERS_43_10_port, B => n2714, S => n1660,
                           Z => n7714);
   U6066 : MUX2_X1 port map( A => REGISTERS_43_9_port, B => n2607, S => n1660, 
                           Z => n7715);
   U6067 : MUX2_X1 port map( A => REGISTERS_43_8_port, B => n2596, S => n1660, 
                           Z => n7716);
   U6068 : MUX2_X1 port map( A => REGISTERS_43_7_port, B => n2585, S => n1661, 
                           Z => n7717);
   U6069 : MUX2_X1 port map( A => REGISTERS_43_6_port, B => n2574, S => n1661, 
                           Z => n7718);
   U6070 : MUX2_X1 port map( A => REGISTERS_43_5_port, B => n2563, S => n1661, 
                           Z => n7719);
   U6071 : MUX2_X1 port map( A => REGISTERS_43_4_port, B => n2552, S => n1661, 
                           Z => n7720);
   U6072 : MUX2_X1 port map( A => REGISTERS_43_3_port, B => n1837, S => n1661, 
                           Z => n7721);
   U6073 : MUX2_X1 port map( A => REGISTERS_43_2_port, B => n1826, S => n1661, 
                           Z => n7722);
   U6074 : MUX2_X1 port map( A => REGISTERS_43_1_port, B => n1815, S => n1661, 
                           Z => n7723);
   U6075 : MUX2_X1 port map( A => REGISTERS_43_0_port, B => n1804, S => n1661, 
                           Z => n7724);
   U6076 : MUX2_X1 port map( A => REGISTERS_42_31_port, B => n2951, S => n1662,
                           Z => n7661);
   U6077 : MUX2_X1 port map( A => REGISTERS_42_30_port, B => n2940, S => n1662,
                           Z => n7662);
   U6078 : MUX2_X1 port map( A => REGISTERS_42_29_port, B => n2929, S => n1662,
                           Z => n7663);
   U6079 : MUX2_X1 port map( A => REGISTERS_42_28_port, B => n2913, S => n1662,
                           Z => n7664);
   U6080 : MUX2_X1 port map( A => REGISTERS_42_27_port, B => n2902, S => n1662,
                           Z => n7665);
   U6081 : MUX2_X1 port map( A => REGISTERS_42_26_port, B => n2890, S => n1662,
                           Z => n7666);
   U6082 : MUX2_X1 port map( A => REGISTERS_42_25_port, B => n2879, S => n1662,
                           Z => n7667);
   U6083 : MUX2_X1 port map( A => REGISTERS_42_24_port, B => n2868, S => n1662,
                           Z => n7668);
   U6084 : MUX2_X1 port map( A => REGISTERS_42_23_port, B => n2857, S => n1662,
                           Z => n7669);
   U6085 : MUX2_X1 port map( A => REGISTERS_42_22_port, B => n2846, S => n1662,
                           Z => n7670);
   U6086 : MUX2_X1 port map( A => REGISTERS_42_21_port, B => n2835, S => n1662,
                           Z => n7671);
   U6087 : MUX2_X1 port map( A => REGISTERS_42_20_port, B => n2824, S => n1662,
                           Z => n7672);
   U6088 : MUX2_X1 port map( A => REGISTERS_42_19_port, B => n2813, S => n1663,
                           Z => n7673);
   U6089 : MUX2_X1 port map( A => REGISTERS_42_18_port, B => n2802, S => n1663,
                           Z => n7674);
   U6090 : MUX2_X1 port map( A => REGISTERS_42_17_port, B => n2791, S => n1663,
                           Z => n7675);
   U6091 : MUX2_X1 port map( A => REGISTERS_42_16_port, B => n2780, S => n1663,
                           Z => n7676);
   U6092 : MUX2_X1 port map( A => REGISTERS_42_15_port, B => n2769, S => n1663,
                           Z => n7677);
   U6093 : MUX2_X1 port map( A => REGISTERS_42_14_port, B => n2758, S => n1663,
                           Z => n7678);
   U6094 : MUX2_X1 port map( A => REGISTERS_42_13_port, B => n2747, S => n1663,
                           Z => n7679);
   U6095 : MUX2_X1 port map( A => REGISTERS_42_12_port, B => n2736, S => n1663,
                           Z => n7680);
   U6096 : MUX2_X1 port map( A => REGISTERS_42_11_port, B => n2725, S => n1663,
                           Z => n7681);
   U6097 : MUX2_X1 port map( A => REGISTERS_42_10_port, B => n2714, S => n1663,
                           Z => n7682);
   U6098 : MUX2_X1 port map( A => REGISTERS_42_9_port, B => n2607, S => n1663, 
                           Z => n7683);
   U6099 : MUX2_X1 port map( A => REGISTERS_42_8_port, B => n2596, S => n1663, 
                           Z => n7684);
   U6100 : MUX2_X1 port map( A => REGISTERS_42_7_port, B => n2585, S => n1664, 
                           Z => n7685);
   U6101 : MUX2_X1 port map( A => REGISTERS_42_6_port, B => n2574, S => n1664, 
                           Z => n7686);
   U6102 : MUX2_X1 port map( A => REGISTERS_42_5_port, B => n2563, S => n1664, 
                           Z => n7687);
   U6103 : MUX2_X1 port map( A => REGISTERS_42_4_port, B => n2552, S => n1664, 
                           Z => n7688);
   U6104 : MUX2_X1 port map( A => REGISTERS_42_3_port, B => n1837, S => n1664, 
                           Z => n7689);
   U6105 : MUX2_X1 port map( A => REGISTERS_42_2_port, B => n1826, S => n1664, 
                           Z => n7690);
   U6106 : MUX2_X1 port map( A => REGISTERS_42_1_port, B => n1815, S => n1664, 
                           Z => n7691);
   U6107 : MUX2_X1 port map( A => REGISTERS_42_0_port, B => n1804, S => n1664, 
                           Z => n7692);
   U6108 : MUX2_X1 port map( A => REGISTERS_41_31_port, B => n2951, S => n1665,
                           Z => n7629);
   U6109 : MUX2_X1 port map( A => REGISTERS_41_30_port, B => n2940, S => n1665,
                           Z => n7630);
   U6110 : MUX2_X1 port map( A => REGISTERS_41_29_port, B => n2929, S => n1665,
                           Z => n7631);
   U6111 : MUX2_X1 port map( A => REGISTERS_41_28_port, B => n2913, S => n1665,
                           Z => n7632);
   U6112 : MUX2_X1 port map( A => REGISTERS_41_27_port, B => n2902, S => n1665,
                           Z => n7633);
   U6113 : MUX2_X1 port map( A => REGISTERS_41_26_port, B => n2890, S => n1665,
                           Z => n7634);
   U6114 : MUX2_X1 port map( A => REGISTERS_41_25_port, B => n2879, S => n1665,
                           Z => n7635);
   U6115 : MUX2_X1 port map( A => REGISTERS_41_24_port, B => n2868, S => n1665,
                           Z => n7636);
   U6116 : MUX2_X1 port map( A => REGISTERS_41_23_port, B => n2857, S => n1665,
                           Z => n7637);
   U6117 : MUX2_X1 port map( A => REGISTERS_41_22_port, B => n2846, S => n1665,
                           Z => n7638);
   U6118 : MUX2_X1 port map( A => REGISTERS_41_21_port, B => n2835, S => n1665,
                           Z => n7639);
   U6119 : MUX2_X1 port map( A => REGISTERS_41_20_port, B => n2824, S => n1665,
                           Z => n7640);
   U6120 : MUX2_X1 port map( A => REGISTERS_41_19_port, B => n2813, S => n1666,
                           Z => n7641);
   U6121 : MUX2_X1 port map( A => REGISTERS_41_18_port, B => n2802, S => n1666,
                           Z => n7642);
   U6122 : MUX2_X1 port map( A => REGISTERS_41_17_port, B => n2791, S => n1666,
                           Z => n7643);
   U6123 : MUX2_X1 port map( A => REGISTERS_41_16_port, B => n2780, S => n1666,
                           Z => n7644);
   U6124 : MUX2_X1 port map( A => REGISTERS_41_15_port, B => n2769, S => n1666,
                           Z => n7645);
   U6125 : MUX2_X1 port map( A => REGISTERS_41_14_port, B => n2758, S => n1666,
                           Z => n7646);
   U6126 : MUX2_X1 port map( A => REGISTERS_41_13_port, B => n2747, S => n1666,
                           Z => n7647);
   U6127 : MUX2_X1 port map( A => REGISTERS_41_12_port, B => n2736, S => n1666,
                           Z => n7648);
   U6128 : MUX2_X1 port map( A => REGISTERS_41_11_port, B => n2725, S => n1666,
                           Z => n7649);
   U6129 : MUX2_X1 port map( A => REGISTERS_41_10_port, B => n2714, S => n1666,
                           Z => n7650);
   U6130 : MUX2_X1 port map( A => REGISTERS_41_9_port, B => n2607, S => n1666, 
                           Z => n7651);
   U6131 : MUX2_X1 port map( A => REGISTERS_41_8_port, B => n2596, S => n1666, 
                           Z => n7652);
   U6132 : MUX2_X1 port map( A => REGISTERS_41_7_port, B => n2585, S => n1667, 
                           Z => n7653);
   U6133 : MUX2_X1 port map( A => REGISTERS_41_6_port, B => n2574, S => n1667, 
                           Z => n7654);
   U6134 : MUX2_X1 port map( A => REGISTERS_41_5_port, B => n2563, S => n1667, 
                           Z => n7655);
   U6135 : MUX2_X1 port map( A => REGISTERS_41_4_port, B => n2552, S => n1667, 
                           Z => n7656);
   U6136 : MUX2_X1 port map( A => REGISTERS_41_3_port, B => n1837, S => n1667, 
                           Z => n7657);
   U6137 : MUX2_X1 port map( A => REGISTERS_41_2_port, B => n1826, S => n1667, 
                           Z => n7658);
   U6138 : MUX2_X1 port map( A => REGISTERS_41_1_port, B => n1815, S => n1667, 
                           Z => n7659);
   U6139 : MUX2_X1 port map( A => REGISTERS_41_0_port, B => n1804, S => n1667, 
                           Z => n7660);
   U6140 : MUX2_X1 port map( A => REGISTERS_40_31_port, B => n2951, S => n1668,
                           Z => n7597);
   U6141 : MUX2_X1 port map( A => REGISTERS_40_30_port, B => n2940, S => n1668,
                           Z => n7598);
   U6142 : MUX2_X1 port map( A => REGISTERS_40_29_port, B => n2929, S => n1668,
                           Z => n7599);
   U6143 : MUX2_X1 port map( A => REGISTERS_40_28_port, B => n2913, S => n1668,
                           Z => n7600);
   U6144 : MUX2_X1 port map( A => REGISTERS_40_27_port, B => n2902, S => n1668,
                           Z => n7601);
   U6145 : MUX2_X1 port map( A => REGISTERS_40_26_port, B => n2890, S => n1668,
                           Z => n7602);
   U6146 : MUX2_X1 port map( A => REGISTERS_40_25_port, B => n2879, S => n1668,
                           Z => n7603);
   U6147 : MUX2_X1 port map( A => REGISTERS_40_24_port, B => n2868, S => n1668,
                           Z => n7604);
   U6148 : MUX2_X1 port map( A => REGISTERS_40_23_port, B => n2857, S => n1668,
                           Z => n7605);
   U6149 : MUX2_X1 port map( A => REGISTERS_40_22_port, B => n2846, S => n1668,
                           Z => n7606);
   U6150 : MUX2_X1 port map( A => REGISTERS_40_21_port, B => n2835, S => n1668,
                           Z => n7607);
   U6151 : MUX2_X1 port map( A => REGISTERS_40_20_port, B => n2824, S => n1668,
                           Z => n7608);
   U6152 : MUX2_X1 port map( A => REGISTERS_40_19_port, B => n2813, S => n1669,
                           Z => n7609);
   U6153 : MUX2_X1 port map( A => REGISTERS_40_18_port, B => n2802, S => n1669,
                           Z => n7610);
   U6154 : MUX2_X1 port map( A => REGISTERS_40_17_port, B => n2791, S => n1669,
                           Z => n7611);
   U6155 : MUX2_X1 port map( A => REGISTERS_40_16_port, B => n2780, S => n1669,
                           Z => n7612);
   U6156 : MUX2_X1 port map( A => REGISTERS_40_15_port, B => n2769, S => n1669,
                           Z => n7613);
   U6157 : MUX2_X1 port map( A => REGISTERS_40_14_port, B => n2758, S => n1669,
                           Z => n7614);
   U6158 : MUX2_X1 port map( A => REGISTERS_40_13_port, B => n2747, S => n1669,
                           Z => n7615);
   U6159 : MUX2_X1 port map( A => REGISTERS_40_12_port, B => n2736, S => n1669,
                           Z => n7616);
   U6160 : MUX2_X1 port map( A => REGISTERS_40_11_port, B => n2725, S => n1669,
                           Z => n7617);
   U6161 : MUX2_X1 port map( A => REGISTERS_40_10_port, B => n2714, S => n1669,
                           Z => n7618);
   U6162 : MUX2_X1 port map( A => REGISTERS_40_9_port, B => n2607, S => n1669, 
                           Z => n7619);
   U6163 : MUX2_X1 port map( A => REGISTERS_40_8_port, B => n2596, S => n1669, 
                           Z => n7620);
   U6164 : MUX2_X1 port map( A => REGISTERS_40_7_port, B => n2585, S => n1670, 
                           Z => n7621);
   U6165 : MUX2_X1 port map( A => REGISTERS_40_6_port, B => n2574, S => n1670, 
                           Z => n7622);
   U6166 : MUX2_X1 port map( A => REGISTERS_40_5_port, B => n2563, S => n1670, 
                           Z => n7623);
   U6167 : MUX2_X1 port map( A => REGISTERS_40_4_port, B => n2552, S => n1670, 
                           Z => n7624);
   U6168 : MUX2_X1 port map( A => REGISTERS_40_3_port, B => n1837, S => n1670, 
                           Z => n7625);
   U6169 : MUX2_X1 port map( A => REGISTERS_40_2_port, B => n1826, S => n1670, 
                           Z => n7626);
   U6170 : MUX2_X1 port map( A => REGISTERS_40_1_port, B => n1815, S => n1670, 
                           Z => n7627);
   U6171 : MUX2_X1 port map( A => REGISTERS_40_0_port, B => n1804, S => n1670, 
                           Z => n7628);
   U6172 : MUX2_X1 port map( A => REGISTERS_39_31_port, B => n2951, S => n1671,
                           Z => n7565);
   U6173 : MUX2_X1 port map( A => REGISTERS_39_30_port, B => n2940, S => n1671,
                           Z => n7566);
   U6174 : MUX2_X1 port map( A => REGISTERS_39_29_port, B => n2929, S => n1671,
                           Z => n7567);
   U6175 : MUX2_X1 port map( A => REGISTERS_39_28_port, B => n2913, S => n1671,
                           Z => n7568);
   U6176 : MUX2_X1 port map( A => REGISTERS_39_27_port, B => n2902, S => n1671,
                           Z => n7569);
   U6177 : MUX2_X1 port map( A => REGISTERS_39_26_port, B => n2890, S => n1671,
                           Z => n7570);
   U6178 : MUX2_X1 port map( A => REGISTERS_39_25_port, B => n2879, S => n1671,
                           Z => n7571);
   U6179 : MUX2_X1 port map( A => REGISTERS_39_24_port, B => n2868, S => n1671,
                           Z => n7572);
   U6180 : MUX2_X1 port map( A => REGISTERS_39_23_port, B => n2857, S => n1671,
                           Z => n7573);
   U6181 : MUX2_X1 port map( A => REGISTERS_39_22_port, B => n2846, S => n1671,
                           Z => n7574);
   U6182 : MUX2_X1 port map( A => REGISTERS_39_21_port, B => n2835, S => n1671,
                           Z => n7575);
   U6183 : MUX2_X1 port map( A => REGISTERS_39_20_port, B => n2824, S => n1671,
                           Z => n7576);
   U6184 : MUX2_X1 port map( A => REGISTERS_39_19_port, B => n2813, S => n1672,
                           Z => n7577);
   U6185 : MUX2_X1 port map( A => REGISTERS_39_18_port, B => n2802, S => n1672,
                           Z => n7578);
   U6186 : MUX2_X1 port map( A => REGISTERS_39_17_port, B => n2791, S => n1672,
                           Z => n7579);
   U6187 : MUX2_X1 port map( A => REGISTERS_39_16_port, B => n2780, S => n1672,
                           Z => n7580);
   U6188 : MUX2_X1 port map( A => REGISTERS_39_15_port, B => n2769, S => n1672,
                           Z => n7581);
   U6189 : MUX2_X1 port map( A => REGISTERS_39_14_port, B => n2758, S => n1672,
                           Z => n7582);
   U6190 : MUX2_X1 port map( A => REGISTERS_39_13_port, B => n2747, S => n1672,
                           Z => n7583);
   U6191 : MUX2_X1 port map( A => REGISTERS_39_12_port, B => n2736, S => n1672,
                           Z => n7584);
   U6192 : MUX2_X1 port map( A => REGISTERS_39_11_port, B => n2725, S => n1672,
                           Z => n7585);
   U6193 : MUX2_X1 port map( A => REGISTERS_39_10_port, B => n2714, S => n1672,
                           Z => n7586);
   U6194 : MUX2_X1 port map( A => REGISTERS_39_9_port, B => n2607, S => n1672, 
                           Z => n7587);
   U6195 : MUX2_X1 port map( A => REGISTERS_39_8_port, B => n2596, S => n1672, 
                           Z => n7588);
   U6196 : MUX2_X1 port map( A => REGISTERS_39_7_port, B => n2585, S => n1673, 
                           Z => n7589);
   U6197 : MUX2_X1 port map( A => REGISTERS_39_6_port, B => n2574, S => n1673, 
                           Z => n7590);
   U6198 : MUX2_X1 port map( A => REGISTERS_39_5_port, B => n2563, S => n1673, 
                           Z => n7591);
   U6199 : MUX2_X1 port map( A => REGISTERS_39_4_port, B => n2552, S => n1673, 
                           Z => n7592);
   U6200 : MUX2_X1 port map( A => REGISTERS_39_3_port, B => n1837, S => n1673, 
                           Z => n7593);
   U6201 : MUX2_X1 port map( A => REGISTERS_39_2_port, B => n1826, S => n1673, 
                           Z => n7594);
   U6202 : MUX2_X1 port map( A => REGISTERS_39_1_port, B => n1815, S => n1673, 
                           Z => n7595);
   U6203 : MUX2_X1 port map( A => REGISTERS_39_0_port, B => n1804, S => n1673, 
                           Z => n7596);
   U6204 : MUX2_X1 port map( A => REGISTERS_38_31_port, B => n2951, S => n1674,
                           Z => n7533);
   U6205 : MUX2_X1 port map( A => REGISTERS_38_30_port, B => n2940, S => n1674,
                           Z => n7534);
   U6206 : MUX2_X1 port map( A => REGISTERS_38_29_port, B => n2929, S => n1674,
                           Z => n7535);
   U6207 : MUX2_X1 port map( A => REGISTERS_38_28_port, B => n2913, S => n1674,
                           Z => n7536);
   U6208 : MUX2_X1 port map( A => REGISTERS_38_27_port, B => n2902, S => n1674,
                           Z => n7537);
   U6209 : MUX2_X1 port map( A => REGISTERS_38_26_port, B => n2890, S => n1674,
                           Z => n7538);
   U6210 : MUX2_X1 port map( A => REGISTERS_38_25_port, B => n2879, S => n1674,
                           Z => n7539);
   U6211 : MUX2_X1 port map( A => REGISTERS_38_24_port, B => n2868, S => n1674,
                           Z => n7540);
   U6212 : MUX2_X1 port map( A => REGISTERS_38_23_port, B => n2857, S => n1674,
                           Z => n7541);
   U6213 : MUX2_X1 port map( A => REGISTERS_38_22_port, B => n2846, S => n1674,
                           Z => n7542);
   U6214 : MUX2_X1 port map( A => REGISTERS_38_21_port, B => n2835, S => n1674,
                           Z => n7543);
   U6215 : MUX2_X1 port map( A => REGISTERS_38_20_port, B => n2824, S => n1674,
                           Z => n7544);
   U6216 : MUX2_X1 port map( A => REGISTERS_38_19_port, B => n2813, S => n1675,
                           Z => n7545);
   U6217 : MUX2_X1 port map( A => REGISTERS_38_18_port, B => n2802, S => n1675,
                           Z => n7546);
   U6218 : MUX2_X1 port map( A => REGISTERS_38_17_port, B => n2791, S => n1675,
                           Z => n7547);
   U6219 : MUX2_X1 port map( A => REGISTERS_38_16_port, B => n2780, S => n1675,
                           Z => n7548);
   U6220 : MUX2_X1 port map( A => REGISTERS_38_15_port, B => n2769, S => n1675,
                           Z => n7549);
   U6221 : MUX2_X1 port map( A => REGISTERS_38_14_port, B => n2758, S => n1675,
                           Z => n7550);
   U6222 : MUX2_X1 port map( A => REGISTERS_38_13_port, B => n2747, S => n1675,
                           Z => n7551);
   U6223 : MUX2_X1 port map( A => REGISTERS_38_12_port, B => n2736, S => n1675,
                           Z => n7552);
   U6224 : MUX2_X1 port map( A => REGISTERS_38_11_port, B => n2725, S => n1675,
                           Z => n7553);
   U6225 : MUX2_X1 port map( A => REGISTERS_38_10_port, B => n2714, S => n1675,
                           Z => n7554);
   U6226 : MUX2_X1 port map( A => REGISTERS_38_9_port, B => n2607, S => n1675, 
                           Z => n7555);
   U6227 : MUX2_X1 port map( A => REGISTERS_38_8_port, B => n2596, S => n1675, 
                           Z => n7556);
   U6228 : MUX2_X1 port map( A => REGISTERS_38_7_port, B => n2585, S => n1676, 
                           Z => n7557);
   U6229 : MUX2_X1 port map( A => REGISTERS_38_6_port, B => n2574, S => n1676, 
                           Z => n7558);
   U6230 : MUX2_X1 port map( A => REGISTERS_38_5_port, B => n2563, S => n1676, 
                           Z => n7559);
   U6231 : MUX2_X1 port map( A => REGISTERS_38_4_port, B => n2552, S => n1676, 
                           Z => n7560);
   U6232 : MUX2_X1 port map( A => REGISTERS_38_3_port, B => n1837, S => n1676, 
                           Z => n7561);
   U6233 : MUX2_X1 port map( A => REGISTERS_38_2_port, B => n1826, S => n1676, 
                           Z => n7562);
   U6234 : MUX2_X1 port map( A => REGISTERS_38_1_port, B => n1815, S => n1676, 
                           Z => n7563);
   U6235 : MUX2_X1 port map( A => REGISTERS_38_0_port, B => n1804, S => n1676, 
                           Z => n7564);
   U6236 : MUX2_X1 port map( A => n9990, B => n2951, S => n1677, Z => n7501);
   U6237 : MUX2_X1 port map( A => n9991, B => n2940, S => n1677, Z => n7502);
   U6238 : MUX2_X1 port map( A => n9992, B => n2929, S => n1677, Z => n7503);
   U6239 : MUX2_X1 port map( A => n9993, B => n2913, S => n1677, Z => n7504);
   U6240 : MUX2_X1 port map( A => n9994, B => n2902, S => n1677, Z => n7505);
   U6241 : MUX2_X1 port map( A => n9995, B => n2890, S => n1677, Z => n7506);
   U6242 : MUX2_X1 port map( A => n9996, B => n2879, S => n1677, Z => n7507);
   U6243 : MUX2_X1 port map( A => n9997, B => n2868, S => n1677, Z => n7508);
   U6244 : MUX2_X1 port map( A => n9998, B => n2857, S => n1677, Z => n7509);
   U6245 : MUX2_X1 port map( A => n9999, B => n2846, S => n1677, Z => n7510);
   U6246 : MUX2_X1 port map( A => n10000, B => n2835, S => n1677, Z => n7511);
   U6247 : MUX2_X1 port map( A => n10001, B => n2824, S => n1677, Z => n7512);
   U6248 : MUX2_X1 port map( A => n10002, B => n2813, S => n1678, Z => n7513);
   U6249 : MUX2_X1 port map( A => n10003, B => n2802, S => n1678, Z => n7514);
   U6250 : MUX2_X1 port map( A => n10004, B => n2791, S => n1678, Z => n7515);
   U6251 : MUX2_X1 port map( A => n10005, B => n2780, S => n1678, Z => n7516);
   U6252 : MUX2_X1 port map( A => n10006, B => n2769, S => n1678, Z => n7517);
   U6253 : MUX2_X1 port map( A => n10007, B => n2758, S => n1678, Z => n7518);
   U6254 : MUX2_X1 port map( A => n10008, B => n2747, S => n1678, Z => n7519);
   U6255 : MUX2_X1 port map( A => n10009, B => n2736, S => n1678, Z => n7520);
   U6256 : MUX2_X1 port map( A => n10010, B => n2725, S => n1678, Z => n7521);
   U6257 : MUX2_X1 port map( A => n10011, B => n2714, S => n1678, Z => n7522);
   U6258 : MUX2_X1 port map( A => n10012, B => n2607, S => n1678, Z => n7523);
   U6259 : MUX2_X1 port map( A => n10013, B => n2596, S => n1678, Z => n7524);
   U6260 : MUX2_X1 port map( A => n10014, B => n2585, S => n1679, Z => n7525);
   U6261 : MUX2_X1 port map( A => n10015, B => n2574, S => n1679, Z => n7526);
   U6262 : MUX2_X1 port map( A => n10016, B => n2563, S => n1679, Z => n7527);
   U6263 : MUX2_X1 port map( A => n10017, B => n2552, S => n1679, Z => n7528);
   U6264 : MUX2_X1 port map( A => n10018, B => n1837, S => n1679, Z => n7529);
   U6265 : MUX2_X1 port map( A => n10019, B => n1826, S => n1679, Z => n7530);
   U6266 : MUX2_X1 port map( A => n10020, B => n1815, S => n1679, Z => n7531);
   U6267 : MUX2_X1 port map( A => n10021, B => n1804, S => n1679, Z => n7532);
   U6268 : MUX2_X1 port map( A => n9958, B => n2951, S => n1680, Z => n7469);
   U6269 : MUX2_X1 port map( A => n9959, B => n2940, S => n1680, Z => n7470);
   U6270 : MUX2_X1 port map( A => n9960, B => n2929, S => n1680, Z => n7471);
   U6271 : MUX2_X1 port map( A => n9961, B => n2913, S => n1680, Z => n7472);
   U6272 : MUX2_X1 port map( A => n9962, B => n2902, S => n1680, Z => n7473);
   U6273 : MUX2_X1 port map( A => n9963, B => n2890, S => n1680, Z => n7474);
   U6274 : MUX2_X1 port map( A => n9964, B => n2879, S => n1680, Z => n7475);
   U6275 : MUX2_X1 port map( A => n9965, B => n2868, S => n1680, Z => n7476);
   U6276 : MUX2_X1 port map( A => n9966, B => n2857, S => n1680, Z => n7477);
   U6277 : MUX2_X1 port map( A => n9967, B => n2846, S => n1680, Z => n7478);
   U6278 : MUX2_X1 port map( A => n9968, B => n2835, S => n1680, Z => n7479);
   U6279 : MUX2_X1 port map( A => n9969, B => n2824, S => n1680, Z => n7480);
   U6280 : MUX2_X1 port map( A => n9970, B => n2813, S => n1681, Z => n7481);
   U6281 : MUX2_X1 port map( A => n9971, B => n2802, S => n1681, Z => n7482);
   U6282 : MUX2_X1 port map( A => n9972, B => n2791, S => n1681, Z => n7483);
   U6283 : MUX2_X1 port map( A => n9973, B => n2780, S => n1681, Z => n7484);
   U6284 : MUX2_X1 port map( A => n9974, B => n2769, S => n1681, Z => n7485);
   U6285 : MUX2_X1 port map( A => n9975, B => n2758, S => n1681, Z => n7486);
   U6286 : MUX2_X1 port map( A => n9976, B => n2747, S => n1681, Z => n7487);
   U6287 : MUX2_X1 port map( A => n9977, B => n2736, S => n1681, Z => n7488);
   U6288 : MUX2_X1 port map( A => n9978, B => n2725, S => n1681, Z => n7489);
   U6289 : MUX2_X1 port map( A => n9979, B => n2714, S => n1681, Z => n7490);
   U6290 : MUX2_X1 port map( A => n9980, B => n2607, S => n1681, Z => n7491);
   U6291 : MUX2_X1 port map( A => n9981, B => n2596, S => n1681, Z => n7492);
   U6292 : MUX2_X1 port map( A => n9982, B => n2585, S => n1682, Z => n7493);
   U6293 : MUX2_X1 port map( A => n9983, B => n2574, S => n1682, Z => n7494);
   U6294 : MUX2_X1 port map( A => n9984, B => n2563, S => n1682, Z => n7495);
   U6295 : MUX2_X1 port map( A => n9985, B => n2552, S => n1682, Z => n7496);
   U6296 : MUX2_X1 port map( A => n9986, B => n1837, S => n1682, Z => n7497);
   U6297 : MUX2_X1 port map( A => n9987, B => n1826, S => n1682, Z => n7498);
   U6298 : MUX2_X1 port map( A => n9988, B => n1815, S => n1682, Z => n7499);
   U6299 : MUX2_X1 port map( A => n9989, B => n1804, S => n1682, Z => n7500);
   U6300 : MUX2_X1 port map( A => n9926, B => n2951, S => n1683, Z => n7437);
   U6301 : MUX2_X1 port map( A => n9927, B => n2940, S => n1683, Z => n7438);
   U6302 : MUX2_X1 port map( A => n9928, B => n2929, S => n1683, Z => n7439);
   U6303 : MUX2_X1 port map( A => n9929, B => n2913, S => n1683, Z => n7440);
   U6304 : MUX2_X1 port map( A => n9930, B => n2902, S => n1683, Z => n7441);
   U6305 : MUX2_X1 port map( A => n9931, B => n2890, S => n1683, Z => n7442);
   U6306 : MUX2_X1 port map( A => n9932, B => n2879, S => n1683, Z => n7443);
   U6307 : MUX2_X1 port map( A => n9933, B => n2868, S => n1683, Z => n7444);
   U6308 : MUX2_X1 port map( A => n9934, B => n2857, S => n1683, Z => n7445);
   U6309 : MUX2_X1 port map( A => n9935, B => n2846, S => n1683, Z => n7446);
   U6310 : MUX2_X1 port map( A => n9936, B => n2835, S => n1683, Z => n7447);
   U6311 : MUX2_X1 port map( A => n9937, B => n2824, S => n1683, Z => n7448);
   U6312 : MUX2_X1 port map( A => n9938, B => n2813, S => n1684, Z => n7449);
   U6313 : MUX2_X1 port map( A => n9939, B => n2802, S => n1684, Z => n7450);
   U6314 : MUX2_X1 port map( A => n9940, B => n2791, S => n1684, Z => n7451);
   U6315 : MUX2_X1 port map( A => n9941, B => n2780, S => n1684, Z => n7452);
   U6316 : MUX2_X1 port map( A => n9942, B => n2769, S => n1684, Z => n7453);
   U6317 : MUX2_X1 port map( A => n9943, B => n2758, S => n1684, Z => n7454);
   U6318 : MUX2_X1 port map( A => n9944, B => n2747, S => n1684, Z => n7455);
   U6319 : MUX2_X1 port map( A => n9945, B => n2736, S => n1684, Z => n7456);
   U6320 : MUX2_X1 port map( A => n9946, B => n2725, S => n1684, Z => n7457);
   U6321 : MUX2_X1 port map( A => n9947, B => n2714, S => n1684, Z => n7458);
   U6322 : MUX2_X1 port map( A => n9948, B => n2607, S => n1684, Z => n7459);
   U6323 : MUX2_X1 port map( A => n9949, B => n2596, S => n1684, Z => n7460);
   U6324 : MUX2_X1 port map( A => n9950, B => n2585, S => n1685, Z => n7461);
   U6325 : MUX2_X1 port map( A => n9951, B => n2574, S => n1685, Z => n7462);
   U6326 : MUX2_X1 port map( A => n9952, B => n2563, S => n1685, Z => n7463);
   U6327 : MUX2_X1 port map( A => n9953, B => n2552, S => n1685, Z => n7464);
   U6328 : MUX2_X1 port map( A => n9954, B => n1837, S => n1685, Z => n7465);
   U6329 : MUX2_X1 port map( A => n9955, B => n1826, S => n1685, Z => n7466);
   U6330 : MUX2_X1 port map( A => n9956, B => n1815, S => n1685, Z => n7467);
   U6331 : MUX2_X1 port map( A => n9957, B => n1804, S => n1685, Z => n7468);
   U6332 : MUX2_X1 port map( A => REGISTERS_34_31_port, B => n2951, S => n1686,
                           Z => n7405);
   U6333 : MUX2_X1 port map( A => REGISTERS_34_30_port, B => n2940, S => n1686,
                           Z => n7406);
   U6334 : MUX2_X1 port map( A => REGISTERS_34_29_port, B => n2929, S => n1686,
                           Z => n7407);
   U6335 : MUX2_X1 port map( A => REGISTERS_34_28_port, B => n2913, S => n1686,
                           Z => n7408);
   U6336 : MUX2_X1 port map( A => REGISTERS_34_27_port, B => n2902, S => n1686,
                           Z => n7409);
   U6337 : MUX2_X1 port map( A => REGISTERS_34_26_port, B => n2890, S => n1686,
                           Z => n7410);
   U6338 : MUX2_X1 port map( A => REGISTERS_34_25_port, B => n2879, S => n1686,
                           Z => n7411);
   U6339 : MUX2_X1 port map( A => REGISTERS_34_24_port, B => n2868, S => n1686,
                           Z => n7412);
   U6340 : MUX2_X1 port map( A => REGISTERS_34_23_port, B => n2857, S => n1686,
                           Z => n7413);
   U6341 : MUX2_X1 port map( A => REGISTERS_34_22_port, B => n2846, S => n1686,
                           Z => n7414);
   U6342 : MUX2_X1 port map( A => REGISTERS_34_21_port, B => n2835, S => n1686,
                           Z => n7415);
   U6343 : MUX2_X1 port map( A => REGISTERS_34_20_port, B => n2824, S => n1686,
                           Z => n7416);
   U6344 : MUX2_X1 port map( A => REGISTERS_34_19_port, B => n2813, S => n1687,
                           Z => n7417);
   U6345 : MUX2_X1 port map( A => REGISTERS_34_18_port, B => n2802, S => n1687,
                           Z => n7418);
   U6346 : MUX2_X1 port map( A => REGISTERS_34_17_port, B => n2791, S => n1687,
                           Z => n7419);
   U6347 : MUX2_X1 port map( A => REGISTERS_34_16_port, B => n2780, S => n1687,
                           Z => n7420);
   U6348 : MUX2_X1 port map( A => REGISTERS_34_15_port, B => n2769, S => n1687,
                           Z => n7421);
   U6349 : MUX2_X1 port map( A => REGISTERS_34_14_port, B => n2758, S => n1687,
                           Z => n7422);
   U6350 : MUX2_X1 port map( A => REGISTERS_34_13_port, B => n2747, S => n1687,
                           Z => n7423);
   U6351 : MUX2_X1 port map( A => REGISTERS_34_12_port, B => n2736, S => n1687,
                           Z => n7424);
   U6352 : MUX2_X1 port map( A => REGISTERS_34_11_port, B => n2725, S => n1687,
                           Z => n7425);
   U6353 : MUX2_X1 port map( A => REGISTERS_34_10_port, B => n2714, S => n1687,
                           Z => n7426);
   U6354 : MUX2_X1 port map( A => REGISTERS_34_9_port, B => n2607, S => n1687, 
                           Z => n7427);
   U6355 : MUX2_X1 port map( A => REGISTERS_34_8_port, B => n2596, S => n1687, 
                           Z => n7428);
   U6356 : MUX2_X1 port map( A => REGISTERS_34_7_port, B => n2585, S => n1688, 
                           Z => n7429);
   U6357 : MUX2_X1 port map( A => REGISTERS_34_6_port, B => n2574, S => n1688, 
                           Z => n7430);
   U6358 : MUX2_X1 port map( A => REGISTERS_34_5_port, B => n2563, S => n1688, 
                           Z => n7431);
   U6359 : MUX2_X1 port map( A => REGISTERS_34_4_port, B => n2552, S => n1688, 
                           Z => n7432);
   U6360 : MUX2_X1 port map( A => REGISTERS_34_3_port, B => n1837, S => n1688, 
                           Z => n7433);
   U6361 : MUX2_X1 port map( A => REGISTERS_34_2_port, B => n1826, S => n1688, 
                           Z => n7434);
   U6362 : MUX2_X1 port map( A => REGISTERS_34_1_port, B => n1815, S => n1688, 
                           Z => n7435);
   U6363 : MUX2_X1 port map( A => REGISTERS_34_0_port, B => n1804, S => n1688, 
                           Z => n7436);
   U6364 : MUX2_X1 port map( A => REGISTERS_33_31_port, B => n2951, S => n1689,
                           Z => n7373);
   U6365 : MUX2_X1 port map( A => REGISTERS_33_30_port, B => n2940, S => n1689,
                           Z => n7374);
   U6366 : MUX2_X1 port map( A => REGISTERS_33_29_port, B => n2929, S => n1689,
                           Z => n7375);
   U6367 : MUX2_X1 port map( A => REGISTERS_33_28_port, B => n2913, S => n1689,
                           Z => n7376);
   U6368 : MUX2_X1 port map( A => REGISTERS_33_27_port, B => n2902, S => n1689,
                           Z => n7377);
   U6369 : MUX2_X1 port map( A => REGISTERS_33_26_port, B => n2890, S => n1689,
                           Z => n7378);
   U6370 : MUX2_X1 port map( A => REGISTERS_33_25_port, B => n2879, S => n1689,
                           Z => n7379);
   U6371 : MUX2_X1 port map( A => REGISTERS_33_24_port, B => n2868, S => n1689,
                           Z => n7380);
   U6372 : MUX2_X1 port map( A => REGISTERS_33_23_port, B => n2857, S => n1689,
                           Z => n7381);
   U6373 : MUX2_X1 port map( A => REGISTERS_33_22_port, B => n2846, S => n1689,
                           Z => n7382);
   U6374 : MUX2_X1 port map( A => REGISTERS_33_21_port, B => n2835, S => n1689,
                           Z => n7383);
   U6375 : MUX2_X1 port map( A => REGISTERS_33_20_port, B => n2824, S => n1689,
                           Z => n7384);
   U6376 : MUX2_X1 port map( A => REGISTERS_33_19_port, B => n2813, S => n1690,
                           Z => n7385);
   U6377 : MUX2_X1 port map( A => REGISTERS_33_18_port, B => n2802, S => n1690,
                           Z => n7386);
   U6378 : MUX2_X1 port map( A => REGISTERS_33_17_port, B => n2791, S => n1690,
                           Z => n7387);
   U6379 : MUX2_X1 port map( A => REGISTERS_33_16_port, B => n2780, S => n1690,
                           Z => n7388);
   U6380 : MUX2_X1 port map( A => REGISTERS_33_15_port, B => n2769, S => n1690,
                           Z => n7389);
   U6381 : MUX2_X1 port map( A => REGISTERS_33_14_port, B => n2758, S => n1690,
                           Z => n7390);
   U6382 : MUX2_X1 port map( A => REGISTERS_33_13_port, B => n2747, S => n1690,
                           Z => n7391);
   U6383 : MUX2_X1 port map( A => REGISTERS_33_12_port, B => n2736, S => n1690,
                           Z => n7392);
   U6384 : MUX2_X1 port map( A => REGISTERS_33_11_port, B => n2725, S => n1690,
                           Z => n7393);
   U6385 : MUX2_X1 port map( A => REGISTERS_33_10_port, B => n2714, S => n1690,
                           Z => n7394);
   U6386 : MUX2_X1 port map( A => REGISTERS_33_9_port, B => n2607, S => n1690, 
                           Z => n7395);
   U6387 : MUX2_X1 port map( A => REGISTERS_33_8_port, B => n2596, S => n1690, 
                           Z => n7396);
   U6388 : MUX2_X1 port map( A => REGISTERS_33_7_port, B => n2585, S => n1691, 
                           Z => n7397);
   U6389 : MUX2_X1 port map( A => REGISTERS_33_6_port, B => n2574, S => n1691, 
                           Z => n7398);
   U6390 : MUX2_X1 port map( A => REGISTERS_33_5_port, B => n2563, S => n1691, 
                           Z => n7399);
   U6391 : MUX2_X1 port map( A => REGISTERS_33_4_port, B => n2552, S => n1691, 
                           Z => n7400);
   U6392 : MUX2_X1 port map( A => REGISTERS_33_3_port, B => n1837, S => n1691, 
                           Z => n7401);
   U6393 : MUX2_X1 port map( A => REGISTERS_33_2_port, B => n1826, S => n1691, 
                           Z => n7402);
   U6394 : MUX2_X1 port map( A => REGISTERS_33_1_port, B => n1815, S => n1691, 
                           Z => n7403);
   U6395 : MUX2_X1 port map( A => REGISTERS_33_0_port, B => n1804, S => n1691, 
                           Z => n7404);
   U6396 : MUX2_X1 port map( A => n9894, B => n2952, S => n1692, Z => n7341);
   U6397 : MUX2_X1 port map( A => n9895, B => n2941, S => n1692, Z => n7342);
   U6398 : MUX2_X1 port map( A => n9896, B => n2930, S => n1692, Z => n7343);
   U6399 : MUX2_X1 port map( A => n9897, B => n2914, S => n1692, Z => n7344);
   U6400 : MUX2_X1 port map( A => n9898, B => n2903, S => n1692, Z => n7345);
   U6401 : MUX2_X1 port map( A => n9899, B => n2891, S => n1692, Z => n7346);
   U6402 : MUX2_X1 port map( A => n9900, B => n2880, S => n1692, Z => n7347);
   U6403 : MUX2_X1 port map( A => n9901, B => n2869, S => n1692, Z => n7348);
   U6404 : MUX2_X1 port map( A => n9902, B => n2858, S => n1692, Z => n7349);
   U6405 : MUX2_X1 port map( A => n9903, B => n2847, S => n1692, Z => n7350);
   U6406 : MUX2_X1 port map( A => n9904, B => n2836, S => n1692, Z => n7351);
   U6407 : MUX2_X1 port map( A => n9905, B => n2825, S => n1692, Z => n7352);
   U6408 : MUX2_X1 port map( A => n9906, B => n2814, S => n1693, Z => n7353);
   U6409 : MUX2_X1 port map( A => n9907, B => n2803, S => n1693, Z => n7354);
   U6410 : MUX2_X1 port map( A => n9908, B => n2792, S => n1693, Z => n7355);
   U6411 : MUX2_X1 port map( A => n9909, B => n2781, S => n1693, Z => n7356);
   U6412 : MUX2_X1 port map( A => n9910, B => n2770, S => n1693, Z => n7357);
   U6413 : MUX2_X1 port map( A => n9911, B => n2759, S => n1693, Z => n7358);
   U6414 : MUX2_X1 port map( A => n9912, B => n2748, S => n1693, Z => n7359);
   U6415 : MUX2_X1 port map( A => n9913, B => n2737, S => n1693, Z => n7360);
   U6416 : MUX2_X1 port map( A => n9914, B => n2726, S => n1693, Z => n7361);
   U6417 : MUX2_X1 port map( A => n9915, B => n2715, S => n1693, Z => n7362);
   U6418 : MUX2_X1 port map( A => n9916, B => n2704, S => n1693, Z => n7363);
   U6419 : MUX2_X1 port map( A => n9917, B => n2597, S => n1693, Z => n7364);
   U6420 : MUX2_X1 port map( A => n9918, B => n2586, S => n1694, Z => n7365);
   U6421 : MUX2_X1 port map( A => n9919, B => n2575, S => n1694, Z => n7366);
   U6422 : MUX2_X1 port map( A => n9920, B => n2564, S => n1694, Z => n7367);
   U6423 : MUX2_X1 port map( A => n9921, B => n2553, S => n1694, Z => n7368);
   U6424 : MUX2_X1 port map( A => n9922, B => n1838, S => n1694, Z => n7369);
   U6425 : MUX2_X1 port map( A => n9923, B => n1827, S => n1694, Z => n7370);
   U6426 : MUX2_X1 port map( A => n9924, B => n1816, S => n1694, Z => n7371);
   U6427 : MUX2_X1 port map( A => n9925, B => n1805, S => n1694, Z => n7372);
   U6428 : MUX2_X1 port map( A => n9862, B => n2952, S => n1695, Z => n7309);
   U6429 : MUX2_X1 port map( A => n9863, B => n2941, S => n1695, Z => n7310);
   U6430 : MUX2_X1 port map( A => n9864, B => n2930, S => n1695, Z => n7311);
   U6431 : MUX2_X1 port map( A => n9865, B => n2914, S => n1695, Z => n7312);
   U6432 : MUX2_X1 port map( A => n9866, B => n2903, S => n1695, Z => n7313);
   U6433 : MUX2_X1 port map( A => n9867, B => n2891, S => n1695, Z => n7314);
   U6434 : MUX2_X1 port map( A => n9868, B => n2880, S => n1695, Z => n7315);
   U6435 : MUX2_X1 port map( A => n9869, B => n2869, S => n1695, Z => n7316);
   U6436 : MUX2_X1 port map( A => n9870, B => n2858, S => n1695, Z => n7317);
   U6437 : MUX2_X1 port map( A => n9871, B => n2847, S => n1695, Z => n7318);
   U6438 : MUX2_X1 port map( A => n9872, B => n2836, S => n1695, Z => n7319);
   U6439 : MUX2_X1 port map( A => n9873, B => n2825, S => n1695, Z => n7320);
   U6440 : MUX2_X1 port map( A => n9874, B => n2814, S => n1696, Z => n7321);
   U6441 : MUX2_X1 port map( A => n9875, B => n2803, S => n1696, Z => n7322);
   U6442 : MUX2_X1 port map( A => n9876, B => n2792, S => n1696, Z => n7323);
   U6443 : MUX2_X1 port map( A => n9877, B => n2781, S => n1696, Z => n7324);
   U6444 : MUX2_X1 port map( A => n9878, B => n2770, S => n1696, Z => n7325);
   U6445 : MUX2_X1 port map( A => n9879, B => n2759, S => n1696, Z => n7326);
   U6446 : MUX2_X1 port map( A => n9880, B => n2748, S => n1696, Z => n7327);
   U6447 : MUX2_X1 port map( A => n9881, B => n2737, S => n1696, Z => n7328);
   U6448 : MUX2_X1 port map( A => n9882, B => n2726, S => n1696, Z => n7329);
   U6449 : MUX2_X1 port map( A => n9883, B => n2715, S => n1696, Z => n7330);
   U6450 : MUX2_X1 port map( A => n9884, B => n2704, S => n1696, Z => n7331);
   U6451 : MUX2_X1 port map( A => n9885, B => n2597, S => n1696, Z => n7332);
   U6452 : MUX2_X1 port map( A => n9886, B => n2586, S => n1697, Z => n7333);
   U6453 : MUX2_X1 port map( A => n9887, B => n2575, S => n1697, Z => n7334);
   U6454 : MUX2_X1 port map( A => n9888, B => n2564, S => n1697, Z => n7335);
   U6455 : MUX2_X1 port map( A => n9889, B => n2553, S => n1697, Z => n7336);
   U6456 : MUX2_X1 port map( A => n9890, B => n1838, S => n1697, Z => n7337);
   U6457 : MUX2_X1 port map( A => n9891, B => n1827, S => n1697, Z => n7338);
   U6458 : MUX2_X1 port map( A => n9892, B => n1816, S => n1697, Z => n7339);
   U6459 : MUX2_X1 port map( A => n9893, B => n1805, S => n1697, Z => n7340);
   U6460 : MUX2_X1 port map( A => n9830, B => n2952, S => n1698, Z => n7277);
   U6461 : MUX2_X1 port map( A => n9831, B => n2941, S => n1698, Z => n7278);
   U6462 : MUX2_X1 port map( A => n9832, B => n2930, S => n1698, Z => n7279);
   U6463 : MUX2_X1 port map( A => n9833, B => n2914, S => n1698, Z => n7280);
   U6464 : MUX2_X1 port map( A => n9834, B => n2903, S => n1698, Z => n7281);
   U6465 : MUX2_X1 port map( A => n9835, B => n2891, S => n1698, Z => n7282);
   U6466 : MUX2_X1 port map( A => n9836, B => n2880, S => n1698, Z => n7283);
   U6467 : MUX2_X1 port map( A => n9837, B => n2869, S => n1698, Z => n7284);
   U6468 : MUX2_X1 port map( A => n9838, B => n2858, S => n1698, Z => n7285);
   U6469 : MUX2_X1 port map( A => n9839, B => n2847, S => n1698, Z => n7286);
   U6470 : MUX2_X1 port map( A => n9840, B => n2836, S => n1698, Z => n7287);
   U6471 : MUX2_X1 port map( A => n9841, B => n2825, S => n1698, Z => n7288);
   U6472 : MUX2_X1 port map( A => n9842, B => n2814, S => n1699, Z => n7289);
   U6473 : MUX2_X1 port map( A => n9843, B => n2803, S => n1699, Z => n7290);
   U6474 : MUX2_X1 port map( A => n9844, B => n2792, S => n1699, Z => n7291);
   U6475 : MUX2_X1 port map( A => n9845, B => n2781, S => n1699, Z => n7292);
   U6476 : MUX2_X1 port map( A => n9846, B => n2770, S => n1699, Z => n7293);
   U6477 : MUX2_X1 port map( A => n9847, B => n2759, S => n1699, Z => n7294);
   U6478 : MUX2_X1 port map( A => n9848, B => n2748, S => n1699, Z => n7295);
   U6479 : MUX2_X1 port map( A => n9849, B => n2737, S => n1699, Z => n7296);
   U6480 : MUX2_X1 port map( A => n9850, B => n2726, S => n1699, Z => n7297);
   U6481 : MUX2_X1 port map( A => n9851, B => n2715, S => n1699, Z => n7298);
   U6482 : MUX2_X1 port map( A => n9852, B => n2704, S => n1699, Z => n7299);
   U6483 : MUX2_X1 port map( A => n9853, B => n2597, S => n1699, Z => n7300);
   U6484 : MUX2_X1 port map( A => n9854, B => n2586, S => n1700, Z => n7301);
   U6485 : MUX2_X1 port map( A => n9855, B => n2575, S => n1700, Z => n7302);
   U6486 : MUX2_X1 port map( A => n9856, B => n2564, S => n1700, Z => n7303);
   U6487 : MUX2_X1 port map( A => n9857, B => n2553, S => n1700, Z => n7304);
   U6488 : MUX2_X1 port map( A => n9858, B => n1838, S => n1700, Z => n7305);
   U6489 : MUX2_X1 port map( A => n9859, B => n1827, S => n1700, Z => n7306);
   U6490 : MUX2_X1 port map( A => n9860, B => n1816, S => n1700, Z => n7307);
   U6491 : MUX2_X1 port map( A => n9861, B => n1805, S => n1700, Z => n7308);
   U6492 : MUX2_X1 port map( A => n9798, B => n2952, S => n1701, Z => n7245);
   U6493 : MUX2_X1 port map( A => n9799, B => n2941, S => n1701, Z => n7246);
   U6494 : MUX2_X1 port map( A => n9800, B => n2930, S => n1701, Z => n7247);
   U6495 : MUX2_X1 port map( A => n9801, B => n2914, S => n1701, Z => n7248);
   U6496 : MUX2_X1 port map( A => n9802, B => n2903, S => n1701, Z => n7249);
   U6497 : MUX2_X1 port map( A => n9803, B => n2891, S => n1701, Z => n7250);
   U6498 : MUX2_X1 port map( A => n9804, B => n2880, S => n1701, Z => n7251);
   U6499 : MUX2_X1 port map( A => n9805, B => n2869, S => n1701, Z => n7252);
   U6500 : MUX2_X1 port map( A => n9806, B => n2858, S => n1701, Z => n7253);
   U6501 : MUX2_X1 port map( A => n9807, B => n2847, S => n1701, Z => n7254);
   U6502 : MUX2_X1 port map( A => n9808, B => n2836, S => n1701, Z => n7255);
   U6503 : MUX2_X1 port map( A => n9809, B => n2825, S => n1701, Z => n7256);
   U6504 : MUX2_X1 port map( A => n9810, B => n2814, S => n1702, Z => n7257);
   U6505 : MUX2_X1 port map( A => n9811, B => n2803, S => n1702, Z => n7258);
   U6506 : MUX2_X1 port map( A => n9812, B => n2792, S => n1702, Z => n7259);
   U6507 : MUX2_X1 port map( A => n9813, B => n2781, S => n1702, Z => n7260);
   U6508 : MUX2_X1 port map( A => n9814, B => n2770, S => n1702, Z => n7261);
   U6509 : MUX2_X1 port map( A => n9815, B => n2759, S => n1702, Z => n7262);
   U6510 : MUX2_X1 port map( A => n9816, B => n2748, S => n1702, Z => n7263);
   U6511 : MUX2_X1 port map( A => n9817, B => n2737, S => n1702, Z => n7264);
   U6512 : MUX2_X1 port map( A => n9818, B => n2726, S => n1702, Z => n7265);
   U6513 : MUX2_X1 port map( A => n9819, B => n2715, S => n1702, Z => n7266);
   U6514 : MUX2_X1 port map( A => n9820, B => n2704, S => n1702, Z => n7267);
   U6515 : MUX2_X1 port map( A => n9821, B => n2597, S => n1702, Z => n7268);
   U6516 : MUX2_X1 port map( A => n9822, B => n2586, S => n1703, Z => n7269);
   U6517 : MUX2_X1 port map( A => n9823, B => n2575, S => n1703, Z => n7270);
   U6518 : MUX2_X1 port map( A => n9824, B => n2564, S => n1703, Z => n7271);
   U6519 : MUX2_X1 port map( A => n9825, B => n2553, S => n1703, Z => n7272);
   U6520 : MUX2_X1 port map( A => n9826, B => n1838, S => n1703, Z => n7273);
   U6521 : MUX2_X1 port map( A => n9827, B => n1827, S => n1703, Z => n7274);
   U6522 : MUX2_X1 port map( A => n9828, B => n1816, S => n1703, Z => n7275);
   U6523 : MUX2_X1 port map( A => n9829, B => n1805, S => n1703, Z => n7276);
   U6524 : MUX2_X1 port map( A => n9766, B => n2952, S => n1704, Z => n7213);
   U6525 : MUX2_X1 port map( A => n9767, B => n2941, S => n1704, Z => n7214);
   U6526 : MUX2_X1 port map( A => n9768, B => n2930, S => n1704, Z => n7215);
   U6527 : MUX2_X1 port map( A => n9769, B => n2914, S => n1704, Z => n7216);
   U6528 : MUX2_X1 port map( A => n9770, B => n2903, S => n1704, Z => n7217);
   U6529 : MUX2_X1 port map( A => n9771, B => n2891, S => n1704, Z => n7218);
   U6530 : MUX2_X1 port map( A => n9772, B => n2880, S => n1704, Z => n7219);
   U6531 : MUX2_X1 port map( A => n9773, B => n2869, S => n1704, Z => n7220);
   U6532 : MUX2_X1 port map( A => n9774, B => n2858, S => n1704, Z => n7221);
   U6533 : MUX2_X1 port map( A => n9775, B => n2847, S => n1704, Z => n7222);
   U6534 : MUX2_X1 port map( A => n9776, B => n2836, S => n1704, Z => n7223);
   U6535 : MUX2_X1 port map( A => n9777, B => n2825, S => n1704, Z => n7224);
   U6536 : MUX2_X1 port map( A => n9778, B => n2814, S => n1705, Z => n7225);
   U6537 : MUX2_X1 port map( A => n9779, B => n2803, S => n1705, Z => n7226);
   U6538 : MUX2_X1 port map( A => n9780, B => n2792, S => n1705, Z => n7227);
   U6539 : MUX2_X1 port map( A => n9781, B => n2781, S => n1705, Z => n7228);
   U6540 : MUX2_X1 port map( A => n9782, B => n2770, S => n1705, Z => n7229);
   U6541 : MUX2_X1 port map( A => n9783, B => n2759, S => n1705, Z => n7230);
   U6542 : MUX2_X1 port map( A => n9784, B => n2748, S => n1705, Z => n7231);
   U6543 : MUX2_X1 port map( A => n9785, B => n2737, S => n1705, Z => n7232);
   U6544 : MUX2_X1 port map( A => n9786, B => n2726, S => n1705, Z => n7233);
   U6545 : MUX2_X1 port map( A => n9787, B => n2715, S => n1705, Z => n7234);
   U6546 : MUX2_X1 port map( A => n9788, B => n2704, S => n1705, Z => n7235);
   U6547 : MUX2_X1 port map( A => n9789, B => n2597, S => n1705, Z => n7236);
   U6548 : MUX2_X1 port map( A => n9790, B => n2586, S => n1706, Z => n7237);
   U6549 : MUX2_X1 port map( A => n9791, B => n2575, S => n1706, Z => n7238);
   U6550 : MUX2_X1 port map( A => n9792, B => n2564, S => n1706, Z => n7239);
   U6551 : MUX2_X1 port map( A => n9793, B => n2553, S => n1706, Z => n7240);
   U6552 : MUX2_X1 port map( A => n9794, B => n1838, S => n1706, Z => n7241);
   U6553 : MUX2_X1 port map( A => n9795, B => n1827, S => n1706, Z => n7242);
   U6554 : MUX2_X1 port map( A => n9796, B => n1816, S => n1706, Z => n7243);
   U6555 : MUX2_X1 port map( A => n9797, B => n1805, S => n1706, Z => n7244);
   U6556 : MUX2_X1 port map( A => n9734, B => n2952, S => n1707, Z => n7181);
   U6557 : MUX2_X1 port map( A => n9735, B => n2941, S => n1707, Z => n7182);
   U6558 : MUX2_X1 port map( A => n9736, B => n2930, S => n1707, Z => n7183);
   U6559 : MUX2_X1 port map( A => n9737, B => n2914, S => n1707, Z => n7184);
   U6560 : MUX2_X1 port map( A => n9738, B => n2903, S => n1707, Z => n7185);
   U6561 : MUX2_X1 port map( A => n9739, B => n2891, S => n1707, Z => n7186);
   U6562 : MUX2_X1 port map( A => n9740, B => n2880, S => n1707, Z => n7187);
   U6563 : MUX2_X1 port map( A => n9741, B => n2869, S => n1707, Z => n7188);
   U6564 : MUX2_X1 port map( A => n9742, B => n2858, S => n1707, Z => n7189);
   U6565 : MUX2_X1 port map( A => n9743, B => n2847, S => n1707, Z => n7190);
   U6566 : MUX2_X1 port map( A => n9744, B => n2836, S => n1707, Z => n7191);
   U6567 : MUX2_X1 port map( A => n9745, B => n2825, S => n1707, Z => n7192);
   U6568 : MUX2_X1 port map( A => n9746, B => n2814, S => n1708, Z => n7193);
   U6569 : MUX2_X1 port map( A => n9747, B => n2803, S => n1708, Z => n7194);
   U6570 : MUX2_X1 port map( A => n9748, B => n2792, S => n1708, Z => n7195);
   U6571 : MUX2_X1 port map( A => n9749, B => n2781, S => n1708, Z => n7196);
   U6572 : MUX2_X1 port map( A => n9750, B => n2770, S => n1708, Z => n7197);
   U6573 : MUX2_X1 port map( A => n9751, B => n2759, S => n1708, Z => n7198);
   U6574 : MUX2_X1 port map( A => n9752, B => n2748, S => n1708, Z => n7199);
   U6575 : MUX2_X1 port map( A => n9753, B => n2737, S => n1708, Z => n7200);
   U6576 : MUX2_X1 port map( A => n9754, B => n2726, S => n1708, Z => n7201);
   U6577 : MUX2_X1 port map( A => n9755, B => n2715, S => n1708, Z => n7202);
   U6578 : MUX2_X1 port map( A => n9756, B => n2704, S => n1708, Z => n7203);
   U6579 : MUX2_X1 port map( A => n9757, B => n2597, S => n1708, Z => n7204);
   U6580 : MUX2_X1 port map( A => n9758, B => n2586, S => n1709, Z => n7205);
   U6581 : MUX2_X1 port map( A => n9759, B => n2575, S => n1709, Z => n7206);
   U6582 : MUX2_X1 port map( A => n9760, B => n2564, S => n1709, Z => n7207);
   U6583 : MUX2_X1 port map( A => n9761, B => n2553, S => n1709, Z => n7208);
   U6584 : MUX2_X1 port map( A => n9762, B => n1838, S => n1709, Z => n7209);
   U6585 : MUX2_X1 port map( A => n9763, B => n1827, S => n1709, Z => n7210);
   U6586 : MUX2_X1 port map( A => n9764, B => n1816, S => n1709, Z => n7211);
   U6587 : MUX2_X1 port map( A => n9765, B => n1805, S => n1709, Z => n7212);
   U6588 : MUX2_X1 port map( A => n9702, B => n2952, S => n1710, Z => n7149);
   U6589 : MUX2_X1 port map( A => n9703, B => n2941, S => n1710, Z => n7150);
   U6590 : MUX2_X1 port map( A => n9704, B => n2930, S => n1710, Z => n7151);
   U6591 : MUX2_X1 port map( A => n9705, B => n2914, S => n1710, Z => n7152);
   U6592 : MUX2_X1 port map( A => n9706, B => n2903, S => n1710, Z => n7153);
   U6593 : MUX2_X1 port map( A => n9707, B => n2891, S => n1710, Z => n7154);
   U6594 : MUX2_X1 port map( A => n9708, B => n2880, S => n1710, Z => n7155);
   U6595 : MUX2_X1 port map( A => n9709, B => n2869, S => n1710, Z => n7156);
   U6596 : MUX2_X1 port map( A => n9710, B => n2858, S => n1710, Z => n7157);
   U6597 : MUX2_X1 port map( A => n9711, B => n2847, S => n1710, Z => n7158);
   U6598 : MUX2_X1 port map( A => n9712, B => n2836, S => n1710, Z => n7159);
   U6599 : MUX2_X1 port map( A => n9713, B => n2825, S => n1710, Z => n7160);
   U6600 : MUX2_X1 port map( A => n9714, B => n2814, S => n1711, Z => n7161);
   U6601 : MUX2_X1 port map( A => n9715, B => n2803, S => n1711, Z => n7162);
   U6602 : MUX2_X1 port map( A => n9716, B => n2792, S => n1711, Z => n7163);
   U6603 : MUX2_X1 port map( A => n9717, B => n2781, S => n1711, Z => n7164);
   U6604 : MUX2_X1 port map( A => n9718, B => n2770, S => n1711, Z => n7165);
   U6605 : MUX2_X1 port map( A => n9719, B => n2759, S => n1711, Z => n7166);
   U6606 : MUX2_X1 port map( A => n9720, B => n2748, S => n1711, Z => n7167);
   U6607 : MUX2_X1 port map( A => n9721, B => n2737, S => n1711, Z => n7168);
   U6608 : MUX2_X1 port map( A => n9722, B => n2726, S => n1711, Z => n7169);
   U6609 : MUX2_X1 port map( A => n9723, B => n2715, S => n1711, Z => n7170);
   U6610 : MUX2_X1 port map( A => n9724, B => n2704, S => n1711, Z => n7171);
   U6611 : MUX2_X1 port map( A => n9725, B => n2597, S => n1711, Z => n7172);
   U6612 : MUX2_X1 port map( A => n9726, B => n2586, S => n1712, Z => n7173);
   U6613 : MUX2_X1 port map( A => n9727, B => n2575, S => n1712, Z => n7174);
   U6614 : MUX2_X1 port map( A => n9728, B => n2564, S => n1712, Z => n7175);
   U6615 : MUX2_X1 port map( A => n9729, B => n2553, S => n1712, Z => n7176);
   U6616 : MUX2_X1 port map( A => n9730, B => n1838, S => n1712, Z => n7177);
   U6617 : MUX2_X1 port map( A => n9731, B => n1827, S => n1712, Z => n7178);
   U6618 : MUX2_X1 port map( A => n9732, B => n1816, S => n1712, Z => n7179);
   U6619 : MUX2_X1 port map( A => n9733, B => n1805, S => n1712, Z => n7180);
   U6620 : MUX2_X1 port map( A => n9670, B => n2952, S => n1713, Z => n7117);
   U6621 : MUX2_X1 port map( A => n9671, B => n2941, S => n1713, Z => n7118);
   U6622 : MUX2_X1 port map( A => n9672, B => n2930, S => n1713, Z => n7119);
   U6623 : MUX2_X1 port map( A => n9673, B => n2914, S => n1713, Z => n7120);
   U6624 : MUX2_X1 port map( A => n9674, B => n2903, S => n1713, Z => n7121);
   U6625 : MUX2_X1 port map( A => n9675, B => n2891, S => n1713, Z => n7122);
   U6626 : MUX2_X1 port map( A => n9676, B => n2880, S => n1713, Z => n7123);
   U6627 : MUX2_X1 port map( A => n9677, B => n2869, S => n1713, Z => n7124);
   U6628 : MUX2_X1 port map( A => n9678, B => n2858, S => n1713, Z => n7125);
   U6629 : MUX2_X1 port map( A => n9679, B => n2847, S => n1713, Z => n7126);
   U6630 : MUX2_X1 port map( A => n9680, B => n2836, S => n1713, Z => n7127);
   U6631 : MUX2_X1 port map( A => n9681, B => n2825, S => n1713, Z => n7128);
   U6632 : MUX2_X1 port map( A => n9682, B => n2814, S => n1714, Z => n7129);
   U6633 : MUX2_X1 port map( A => n9683, B => n2803, S => n1714, Z => n7130);
   U6634 : MUX2_X1 port map( A => n9684, B => n2792, S => n1714, Z => n7131);
   U6635 : MUX2_X1 port map( A => n9685, B => n2781, S => n1714, Z => n7132);
   U6636 : MUX2_X1 port map( A => n9686, B => n2770, S => n1714, Z => n7133);
   U6637 : MUX2_X1 port map( A => n9687, B => n2759, S => n1714, Z => n7134);
   U6638 : MUX2_X1 port map( A => n9688, B => n2748, S => n1714, Z => n7135);
   U6639 : MUX2_X1 port map( A => n9689, B => n2737, S => n1714, Z => n7136);
   U6640 : MUX2_X1 port map( A => n9690, B => n2726, S => n1714, Z => n7137);
   U6641 : MUX2_X1 port map( A => n9691, B => n2715, S => n1714, Z => n7138);
   U6642 : MUX2_X1 port map( A => n9692, B => n2704, S => n1714, Z => n7139);
   U6643 : MUX2_X1 port map( A => n9693, B => n2597, S => n1714, Z => n7140);
   U6644 : MUX2_X1 port map( A => n9694, B => n2586, S => n1715, Z => n7141);
   U6645 : MUX2_X1 port map( A => n9695, B => n2575, S => n1715, Z => n7142);
   U6646 : MUX2_X1 port map( A => n9696, B => n2564, S => n1715, Z => n7143);
   U6647 : MUX2_X1 port map( A => n9697, B => n2553, S => n1715, Z => n7144);
   U6648 : MUX2_X1 port map( A => n9698, B => n1838, S => n1715, Z => n7145);
   U6649 : MUX2_X1 port map( A => n9699, B => n1827, S => n1715, Z => n7146);
   U6650 : MUX2_X1 port map( A => n9700, B => n1816, S => n1715, Z => n7147);
   U6651 : MUX2_X1 port map( A => n9701, B => n1805, S => n1715, Z => n7148);
   U6652 : MUX2_X1 port map( A => n9638, B => n2952, S => n1716, Z => n7085);
   U6653 : MUX2_X1 port map( A => n9639, B => n2941, S => n1716, Z => n7086);
   U6654 : MUX2_X1 port map( A => n9640, B => n2930, S => n1716, Z => n7087);
   U6655 : MUX2_X1 port map( A => n9641, B => n2914, S => n1716, Z => n7088);
   U6656 : MUX2_X1 port map( A => n9642, B => n2903, S => n1716, Z => n7089);
   U6657 : MUX2_X1 port map( A => n9643, B => n2891, S => n1716, Z => n7090);
   U6658 : MUX2_X1 port map( A => n9644, B => n2880, S => n1716, Z => n7091);
   U6659 : MUX2_X1 port map( A => n9645, B => n2869, S => n1716, Z => n7092);
   U6660 : MUX2_X1 port map( A => n9646, B => n2858, S => n1716, Z => n7093);
   U6661 : MUX2_X1 port map( A => n9647, B => n2847, S => n1716, Z => n7094);
   U6662 : MUX2_X1 port map( A => n9648, B => n2836, S => n1716, Z => n7095);
   U6663 : MUX2_X1 port map( A => n9649, B => n2825, S => n1716, Z => n7096);
   U6664 : MUX2_X1 port map( A => n9650, B => n2814, S => n1717, Z => n7097);
   U6665 : MUX2_X1 port map( A => n9651, B => n2803, S => n1717, Z => n7098);
   U6666 : MUX2_X1 port map( A => n9652, B => n2792, S => n1717, Z => n7099);
   U6667 : MUX2_X1 port map( A => n9653, B => n2781, S => n1717, Z => n7100);
   U6668 : MUX2_X1 port map( A => n9654, B => n2770, S => n1717, Z => n7101);
   U6669 : MUX2_X1 port map( A => n9655, B => n2759, S => n1717, Z => n7102);
   U6670 : MUX2_X1 port map( A => n9656, B => n2748, S => n1717, Z => n7103);
   U6671 : MUX2_X1 port map( A => n9657, B => n2737, S => n1717, Z => n7104);
   U6672 : MUX2_X1 port map( A => n9658, B => n2726, S => n1717, Z => n7105);
   U6673 : MUX2_X1 port map( A => n9659, B => n2715, S => n1717, Z => n7106);
   U6674 : MUX2_X1 port map( A => n9660, B => n2704, S => n1717, Z => n7107);
   U6675 : MUX2_X1 port map( A => n9661, B => n2597, S => n1717, Z => n7108);
   U6676 : MUX2_X1 port map( A => n9662, B => n2586, S => n1718, Z => n7109);
   U6677 : MUX2_X1 port map( A => n9663, B => n2575, S => n1718, Z => n7110);
   U6678 : MUX2_X1 port map( A => n9664, B => n2564, S => n1718, Z => n7111);
   U6679 : MUX2_X1 port map( A => n9665, B => n2553, S => n1718, Z => n7112);
   U6680 : MUX2_X1 port map( A => n9666, B => n1838, S => n1718, Z => n7113);
   U6681 : MUX2_X1 port map( A => n9667, B => n1827, S => n1718, Z => n7114);
   U6682 : MUX2_X1 port map( A => n9668, B => n1816, S => n1718, Z => n7115);
   U6683 : MUX2_X1 port map( A => n9669, B => n1805, S => n1718, Z => n7116);
   U6684 : MUX2_X1 port map( A => n9606, B => n2952, S => n1719, Z => n7053);
   U6685 : MUX2_X1 port map( A => n9607, B => n2941, S => n1719, Z => n7054);
   U6686 : MUX2_X1 port map( A => n9608, B => n2930, S => n1719, Z => n7055);
   U6687 : MUX2_X1 port map( A => n9609, B => n2914, S => n1719, Z => n7056);
   U6688 : MUX2_X1 port map( A => n9610, B => n2903, S => n1719, Z => n7057);
   U6689 : MUX2_X1 port map( A => n9611, B => n2891, S => n1719, Z => n7058);
   U6690 : MUX2_X1 port map( A => n9612, B => n2880, S => n1719, Z => n7059);
   U6691 : MUX2_X1 port map( A => n9613, B => n2869, S => n1719, Z => n7060);
   U6692 : MUX2_X1 port map( A => n9614, B => n2858, S => n1719, Z => n7061);
   U6693 : MUX2_X1 port map( A => n9615, B => n2847, S => n1719, Z => n7062);
   U6694 : MUX2_X1 port map( A => n9616, B => n2836, S => n1719, Z => n7063);
   U6695 : MUX2_X1 port map( A => n9617, B => n2825, S => n1719, Z => n7064);
   U6696 : MUX2_X1 port map( A => n9618, B => n2814, S => n1720, Z => n7065);
   U6697 : MUX2_X1 port map( A => n9619, B => n2803, S => n1720, Z => n7066);
   U6698 : MUX2_X1 port map( A => n9620, B => n2792, S => n1720, Z => n7067);
   U6699 : MUX2_X1 port map( A => n9621, B => n2781, S => n1720, Z => n7068);
   U6700 : MUX2_X1 port map( A => n9622, B => n2770, S => n1720, Z => n7069);
   U6701 : MUX2_X1 port map( A => n9623, B => n2759, S => n1720, Z => n7070);
   U6702 : MUX2_X1 port map( A => n9624, B => n2748, S => n1720, Z => n7071);
   U6703 : MUX2_X1 port map( A => n9625, B => n2737, S => n1720, Z => n7072);
   U6704 : MUX2_X1 port map( A => n9626, B => n2726, S => n1720, Z => n7073);
   U6705 : MUX2_X1 port map( A => n9627, B => n2715, S => n1720, Z => n7074);
   U6706 : MUX2_X1 port map( A => n9628, B => n2704, S => n1720, Z => n7075);
   U6707 : MUX2_X1 port map( A => n9629, B => n2597, S => n1720, Z => n7076);
   U6708 : MUX2_X1 port map( A => n9630, B => n2586, S => n1721, Z => n7077);
   U6709 : MUX2_X1 port map( A => n9631, B => n2575, S => n1721, Z => n7078);
   U6710 : MUX2_X1 port map( A => n9632, B => n2564, S => n1721, Z => n7079);
   U6711 : MUX2_X1 port map( A => n9633, B => n2553, S => n1721, Z => n7080);
   U6712 : MUX2_X1 port map( A => n9634, B => n1838, S => n1721, Z => n7081);
   U6713 : MUX2_X1 port map( A => n9635, B => n1827, S => n1721, Z => n7082);
   U6714 : MUX2_X1 port map( A => n9636, B => n1816, S => n1721, Z => n7083);
   U6715 : MUX2_X1 port map( A => n9637, B => n1805, S => n1721, Z => n7084);
   U6716 : MUX2_X1 port map( A => n9574, B => n2952, S => n1722, Z => n7021);
   U6717 : MUX2_X1 port map( A => n9575, B => n2941, S => n1722, Z => n7022);
   U6718 : MUX2_X1 port map( A => n9576, B => n2930, S => n1722, Z => n7023);
   U6719 : MUX2_X1 port map( A => n9577, B => n2914, S => n1722, Z => n7024);
   U6720 : MUX2_X1 port map( A => n9578, B => n2903, S => n1722, Z => n7025);
   U6721 : MUX2_X1 port map( A => n9579, B => n2891, S => n1722, Z => n7026);
   U6722 : MUX2_X1 port map( A => n9580, B => n2880, S => n1722, Z => n7027);
   U6723 : MUX2_X1 port map( A => n9581, B => n2869, S => n1722, Z => n7028);
   U6724 : MUX2_X1 port map( A => n9582, B => n2858, S => n1722, Z => n7029);
   U6725 : MUX2_X1 port map( A => n9583, B => n2847, S => n1722, Z => n7030);
   U6726 : MUX2_X1 port map( A => n9584, B => n2836, S => n1722, Z => n7031);
   U6727 : MUX2_X1 port map( A => n9585, B => n2825, S => n1722, Z => n7032);
   U6728 : MUX2_X1 port map( A => n9586, B => n2814, S => n1723, Z => n7033);
   U6729 : MUX2_X1 port map( A => n9587, B => n2803, S => n1723, Z => n7034);
   U6730 : MUX2_X1 port map( A => n9588, B => n2792, S => n1723, Z => n7035);
   U6731 : MUX2_X1 port map( A => n9589, B => n2781, S => n1723, Z => n7036);
   U6732 : MUX2_X1 port map( A => n9590, B => n2770, S => n1723, Z => n7037);
   U6733 : MUX2_X1 port map( A => n9591, B => n2759, S => n1723, Z => n7038);
   U6734 : MUX2_X1 port map( A => n9592, B => n2748, S => n1723, Z => n7039);
   U6735 : MUX2_X1 port map( A => n9593, B => n2737, S => n1723, Z => n7040);
   U6736 : MUX2_X1 port map( A => n9594, B => n2726, S => n1723, Z => n7041);
   U6737 : MUX2_X1 port map( A => n9595, B => n2715, S => n1723, Z => n7042);
   U6738 : MUX2_X1 port map( A => n9596, B => n2704, S => n1723, Z => n7043);
   U6739 : MUX2_X1 port map( A => n9597, B => n2597, S => n1723, Z => n7044);
   U6740 : MUX2_X1 port map( A => n9598, B => n2586, S => n1724, Z => n7045);
   U6741 : MUX2_X1 port map( A => n9599, B => n2575, S => n1724, Z => n7046);
   U6742 : MUX2_X1 port map( A => n9600, B => n2564, S => n1724, Z => n7047);
   U6743 : MUX2_X1 port map( A => n9601, B => n2553, S => n1724, Z => n7048);
   U6744 : MUX2_X1 port map( A => n9602, B => n1838, S => n1724, Z => n7049);
   U6745 : MUX2_X1 port map( A => n9603, B => n1827, S => n1724, Z => n7050);
   U6746 : MUX2_X1 port map( A => n9604, B => n1816, S => n1724, Z => n7051);
   U6747 : MUX2_X1 port map( A => n9605, B => n1805, S => n1724, Z => n7052);
   U6748 : MUX2_X1 port map( A => REGISTERS_21_31_port, B => n2953, S => n1725,
                           Z => n6989);
   U6749 : MUX2_X1 port map( A => REGISTERS_21_30_port, B => n2942, S => n1725,
                           Z => n6990);
   U6750 : MUX2_X1 port map( A => REGISTERS_21_29_port, B => n2931, S => n1725,
                           Z => n6991);
   U6751 : MUX2_X1 port map( A => REGISTERS_21_28_port, B => n2915, S => n1725,
                           Z => n6992);
   U6752 : MUX2_X1 port map( A => REGISTERS_21_27_port, B => n2904, S => n1725,
                           Z => n6993);
   U6753 : MUX2_X1 port map( A => REGISTERS_21_26_port, B => n2892, S => n1725,
                           Z => n6994);
   U6754 : MUX2_X1 port map( A => REGISTERS_21_25_port, B => n2881, S => n1725,
                           Z => n6995);
   U6755 : MUX2_X1 port map( A => REGISTERS_21_24_port, B => n2870, S => n1725,
                           Z => n6996);
   U6756 : MUX2_X1 port map( A => REGISTERS_21_23_port, B => n2859, S => n1725,
                           Z => n6997);
   U6757 : MUX2_X1 port map( A => REGISTERS_21_22_port, B => n2848, S => n1725,
                           Z => n6998);
   U6758 : MUX2_X1 port map( A => REGISTERS_21_21_port, B => n2837, S => n1725,
                           Z => n6999);
   U6759 : MUX2_X1 port map( A => REGISTERS_21_20_port, B => n2826, S => n1725,
                           Z => n7000);
   U6760 : MUX2_X1 port map( A => REGISTERS_21_19_port, B => n2815, S => n1726,
                           Z => n7001);
   U6761 : MUX2_X1 port map( A => REGISTERS_21_18_port, B => n2804, S => n1726,
                           Z => n7002);
   U6762 : MUX2_X1 port map( A => REGISTERS_21_17_port, B => n2793, S => n1726,
                           Z => n7003);
   U6763 : MUX2_X1 port map( A => REGISTERS_21_16_port, B => n2782, S => n1726,
                           Z => n7004);
   U6764 : MUX2_X1 port map( A => REGISTERS_21_15_port, B => n2771, S => n1726,
                           Z => n7005);
   U6765 : MUX2_X1 port map( A => REGISTERS_21_14_port, B => n2760, S => n1726,
                           Z => n7006);
   U6766 : MUX2_X1 port map( A => REGISTERS_21_13_port, B => n2749, S => n1726,
                           Z => n7007);
   U6767 : MUX2_X1 port map( A => REGISTERS_21_12_port, B => n2738, S => n1726,
                           Z => n7008);
   U6768 : MUX2_X1 port map( A => REGISTERS_21_11_port, B => n2727, S => n1726,
                           Z => n7009);
   U6769 : MUX2_X1 port map( A => REGISTERS_21_10_port, B => n2716, S => n1726,
                           Z => n7010);
   U6770 : MUX2_X1 port map( A => REGISTERS_21_9_port, B => n2705, S => n1726, 
                           Z => n7011);
   U6771 : MUX2_X1 port map( A => REGISTERS_21_8_port, B => n2598, S => n1726, 
                           Z => n7012);
   U6772 : MUX2_X1 port map( A => REGISTERS_21_7_port, B => n2587, S => n1727, 
                           Z => n7013);
   U6773 : MUX2_X1 port map( A => REGISTERS_21_6_port, B => n2576, S => n1727, 
                           Z => n7014);
   U6774 : MUX2_X1 port map( A => REGISTERS_21_5_port, B => n2565, S => n1727, 
                           Z => n7015);
   U6775 : MUX2_X1 port map( A => REGISTERS_21_4_port, B => n2554, S => n1727, 
                           Z => n7016);
   U6776 : MUX2_X1 port map( A => REGISTERS_21_3_port, B => n1839, S => n1727, 
                           Z => n7017);
   U6777 : MUX2_X1 port map( A => REGISTERS_21_2_port, B => n1828, S => n1727, 
                           Z => n7018);
   U6778 : MUX2_X1 port map( A => REGISTERS_21_1_port, B => n1817, S => n1727, 
                           Z => n7019);
   U6779 : MUX2_X1 port map( A => REGISTERS_21_0_port, B => n1806, S => n1727, 
                           Z => n7020);
   U6780 : MUX2_X1 port map( A => REGISTERS_20_31_port, B => n2953, S => n1728,
                           Z => n6957);
   U6781 : MUX2_X1 port map( A => REGISTERS_20_30_port, B => n2942, S => n1728,
                           Z => n6958);
   U6782 : MUX2_X1 port map( A => REGISTERS_20_29_port, B => n2931, S => n1728,
                           Z => n6959);
   U6783 : MUX2_X1 port map( A => REGISTERS_20_28_port, B => n2915, S => n1728,
                           Z => n6960);
   U6784 : MUX2_X1 port map( A => REGISTERS_20_27_port, B => n2904, S => n1728,
                           Z => n6961);
   U6785 : MUX2_X1 port map( A => REGISTERS_20_26_port, B => n2892, S => n1728,
                           Z => n6962);
   U6786 : MUX2_X1 port map( A => REGISTERS_20_25_port, B => n2881, S => n1728,
                           Z => n6963);
   U6787 : MUX2_X1 port map( A => REGISTERS_20_24_port, B => n2870, S => n1728,
                           Z => n6964);
   U6788 : MUX2_X1 port map( A => REGISTERS_20_23_port, B => n2859, S => n1728,
                           Z => n6965);
   U6789 : MUX2_X1 port map( A => REGISTERS_20_22_port, B => n2848, S => n1728,
                           Z => n6966);
   U6790 : MUX2_X1 port map( A => REGISTERS_20_21_port, B => n2837, S => n1728,
                           Z => n6967);
   U6791 : MUX2_X1 port map( A => REGISTERS_20_20_port, B => n2826, S => n1728,
                           Z => n6968);
   U6792 : MUX2_X1 port map( A => REGISTERS_20_19_port, B => n2815, S => n1729,
                           Z => n6969);
   U6793 : MUX2_X1 port map( A => REGISTERS_20_18_port, B => n2804, S => n1729,
                           Z => n6970);
   U6794 : MUX2_X1 port map( A => REGISTERS_20_17_port, B => n2793, S => n1729,
                           Z => n6971);
   U6795 : MUX2_X1 port map( A => REGISTERS_20_16_port, B => n2782, S => n1729,
                           Z => n6972);
   U6796 : MUX2_X1 port map( A => REGISTERS_20_15_port, B => n2771, S => n1729,
                           Z => n6973);
   U6797 : MUX2_X1 port map( A => REGISTERS_20_14_port, B => n2760, S => n1729,
                           Z => n6974);
   U6798 : MUX2_X1 port map( A => REGISTERS_20_13_port, B => n2749, S => n1729,
                           Z => n6975);
   U6799 : MUX2_X1 port map( A => REGISTERS_20_12_port, B => n2738, S => n1729,
                           Z => n6976);
   U6800 : MUX2_X1 port map( A => REGISTERS_20_11_port, B => n2727, S => n1729,
                           Z => n6977);
   U6801 : MUX2_X1 port map( A => REGISTERS_20_10_port, B => n2716, S => n1729,
                           Z => n6978);
   U6802 : MUX2_X1 port map( A => REGISTERS_20_9_port, B => n2705, S => n1729, 
                           Z => n6979);
   U6803 : MUX2_X1 port map( A => REGISTERS_20_8_port, B => n2598, S => n1729, 
                           Z => n6980);
   U6804 : MUX2_X1 port map( A => REGISTERS_20_7_port, B => n2587, S => n1730, 
                           Z => n6981);
   U6805 : MUX2_X1 port map( A => REGISTERS_20_6_port, B => n2576, S => n1730, 
                           Z => n6982);
   U6806 : MUX2_X1 port map( A => REGISTERS_20_5_port, B => n2565, S => n1730, 
                           Z => n6983);
   U6807 : MUX2_X1 port map( A => REGISTERS_20_4_port, B => n2554, S => n1730, 
                           Z => n6984);
   U6808 : MUX2_X1 port map( A => REGISTERS_20_3_port, B => n1839, S => n1730, 
                           Z => n6985);
   U6809 : MUX2_X1 port map( A => REGISTERS_20_2_port, B => n1828, S => n1730, 
                           Z => n6986);
   U6810 : MUX2_X1 port map( A => REGISTERS_20_1_port, B => n1817, S => n1730, 
                           Z => n6987);
   U6811 : MUX2_X1 port map( A => REGISTERS_20_0_port, B => n1806, S => n1730, 
                           Z => n6988);
   U6812 : MUX2_X1 port map( A => REGISTERS_19_31_port, B => n2953, S => n1731,
                           Z => n6925);
   U6813 : MUX2_X1 port map( A => REGISTERS_19_30_port, B => n2942, S => n1731,
                           Z => n6926);
   U6814 : MUX2_X1 port map( A => REGISTERS_19_29_port, B => n2931, S => n1731,
                           Z => n6927);
   U6815 : MUX2_X1 port map( A => REGISTERS_19_28_port, B => n2915, S => n1731,
                           Z => n6928);
   U6816 : MUX2_X1 port map( A => REGISTERS_19_27_port, B => n2904, S => n1731,
                           Z => n6929);
   U6817 : MUX2_X1 port map( A => REGISTERS_19_26_port, B => n2892, S => n1731,
                           Z => n6930);
   U6818 : MUX2_X1 port map( A => REGISTERS_19_25_port, B => n2881, S => n1731,
                           Z => n6931);
   U6819 : MUX2_X1 port map( A => REGISTERS_19_24_port, B => n2870, S => n1731,
                           Z => n6932);
   U6820 : MUX2_X1 port map( A => REGISTERS_19_23_port, B => n2859, S => n1731,
                           Z => n6933);
   U6821 : MUX2_X1 port map( A => REGISTERS_19_22_port, B => n2848, S => n1731,
                           Z => n6934);
   U6822 : MUX2_X1 port map( A => REGISTERS_19_21_port, B => n2837, S => n1731,
                           Z => n6935);
   U6823 : MUX2_X1 port map( A => REGISTERS_19_20_port, B => n2826, S => n1731,
                           Z => n6936);
   U6824 : MUX2_X1 port map( A => REGISTERS_19_19_port, B => n2815, S => n1732,
                           Z => n6937);
   U6825 : MUX2_X1 port map( A => REGISTERS_19_18_port, B => n2804, S => n1732,
                           Z => n6938);
   U6826 : MUX2_X1 port map( A => REGISTERS_19_17_port, B => n2793, S => n1732,
                           Z => n6939);
   U6827 : MUX2_X1 port map( A => REGISTERS_19_16_port, B => n2782, S => n1732,
                           Z => n6940);
   U6828 : MUX2_X1 port map( A => REGISTERS_19_15_port, B => n2771, S => n1732,
                           Z => n6941);
   U6829 : MUX2_X1 port map( A => REGISTERS_19_14_port, B => n2760, S => n1732,
                           Z => n6942);
   U6830 : MUX2_X1 port map( A => REGISTERS_19_13_port, B => n2749, S => n1732,
                           Z => n6943);
   U6831 : MUX2_X1 port map( A => REGISTERS_19_12_port, B => n2738, S => n1732,
                           Z => n6944);
   U6832 : MUX2_X1 port map( A => REGISTERS_19_11_port, B => n2727, S => n1732,
                           Z => n6945);
   U6833 : MUX2_X1 port map( A => REGISTERS_19_10_port, B => n2716, S => n1732,
                           Z => n6946);
   U6834 : MUX2_X1 port map( A => REGISTERS_19_9_port, B => n2705, S => n1732, 
                           Z => n6947);
   U6835 : MUX2_X1 port map( A => REGISTERS_19_8_port, B => n2598, S => n1732, 
                           Z => n6948);
   U6836 : MUX2_X1 port map( A => REGISTERS_19_7_port, B => n2587, S => n1733, 
                           Z => n6949);
   U6837 : MUX2_X1 port map( A => REGISTERS_19_6_port, B => n2576, S => n1733, 
                           Z => n6950);
   U6838 : MUX2_X1 port map( A => REGISTERS_19_5_port, B => n2565, S => n1733, 
                           Z => n6951);
   U6839 : MUX2_X1 port map( A => REGISTERS_19_4_port, B => n2554, S => n1733, 
                           Z => n6952);
   U6840 : MUX2_X1 port map( A => REGISTERS_19_3_port, B => n1839, S => n1733, 
                           Z => n6953);
   U6841 : MUX2_X1 port map( A => REGISTERS_19_2_port, B => n1828, S => n1733, 
                           Z => n6954);
   U6842 : MUX2_X1 port map( A => REGISTERS_19_1_port, B => n1817, S => n1733, 
                           Z => n6955);
   U6843 : MUX2_X1 port map( A => REGISTERS_19_0_port, B => n1806, S => n1733, 
                           Z => n6956);
   U6844 : MUX2_X1 port map( A => REGISTERS_18_31_port, B => n2953, S => n1734,
                           Z => n6893);
   U6845 : MUX2_X1 port map( A => REGISTERS_18_30_port, B => n2942, S => n1734,
                           Z => n6894);
   U6846 : MUX2_X1 port map( A => REGISTERS_18_29_port, B => n2931, S => n1734,
                           Z => n6895);
   U6847 : MUX2_X1 port map( A => REGISTERS_18_28_port, B => n2915, S => n1734,
                           Z => n6896);
   U6848 : MUX2_X1 port map( A => REGISTERS_18_27_port, B => n2904, S => n1734,
                           Z => n6897);
   U6849 : MUX2_X1 port map( A => REGISTERS_18_26_port, B => n2892, S => n1734,
                           Z => n6898);
   U6850 : MUX2_X1 port map( A => REGISTERS_18_25_port, B => n2881, S => n1734,
                           Z => n6899);
   U6851 : MUX2_X1 port map( A => REGISTERS_18_24_port, B => n2870, S => n1734,
                           Z => n6900);
   U6852 : MUX2_X1 port map( A => REGISTERS_18_23_port, B => n2859, S => n1734,
                           Z => n6901);
   U6853 : MUX2_X1 port map( A => REGISTERS_18_22_port, B => n2848, S => n1734,
                           Z => n6902);
   U6854 : MUX2_X1 port map( A => REGISTERS_18_21_port, B => n2837, S => n1734,
                           Z => n6903);
   U6855 : MUX2_X1 port map( A => REGISTERS_18_20_port, B => n2826, S => n1734,
                           Z => n6904);
   U6856 : MUX2_X1 port map( A => REGISTERS_18_19_port, B => n2815, S => n1735,
                           Z => n6905);
   U6857 : MUX2_X1 port map( A => REGISTERS_18_18_port, B => n2804, S => n1735,
                           Z => n6906);
   U6858 : MUX2_X1 port map( A => REGISTERS_18_17_port, B => n2793, S => n1735,
                           Z => n6907);
   U6859 : MUX2_X1 port map( A => REGISTERS_18_16_port, B => n2782, S => n1735,
                           Z => n6908);
   U6860 : MUX2_X1 port map( A => REGISTERS_18_15_port, B => n2771, S => n1735,
                           Z => n6909);
   U6861 : MUX2_X1 port map( A => REGISTERS_18_14_port, B => n2760, S => n1735,
                           Z => n6910);
   U6862 : MUX2_X1 port map( A => REGISTERS_18_13_port, B => n2749, S => n1735,
                           Z => n6911);
   U6863 : MUX2_X1 port map( A => REGISTERS_18_12_port, B => n2738, S => n1735,
                           Z => n6912);
   U6864 : MUX2_X1 port map( A => REGISTERS_18_11_port, B => n2727, S => n1735,
                           Z => n6913);
   U6865 : MUX2_X1 port map( A => REGISTERS_18_10_port, B => n2716, S => n1735,
                           Z => n6914);
   U6866 : MUX2_X1 port map( A => REGISTERS_18_9_port, B => n2705, S => n1735, 
                           Z => n6915);
   U6867 : MUX2_X1 port map( A => REGISTERS_18_8_port, B => n2598, S => n1735, 
                           Z => n6916);
   U6868 : MUX2_X1 port map( A => REGISTERS_18_7_port, B => n2587, S => n1736, 
                           Z => n6917);
   U6869 : MUX2_X1 port map( A => REGISTERS_18_6_port, B => n2576, S => n1736, 
                           Z => n6918);
   U6870 : MUX2_X1 port map( A => REGISTERS_18_5_port, B => n2565, S => n1736, 
                           Z => n6919);
   U6871 : MUX2_X1 port map( A => REGISTERS_18_4_port, B => n2554, S => n1736, 
                           Z => n6920);
   U6872 : MUX2_X1 port map( A => REGISTERS_18_3_port, B => n1839, S => n1736, 
                           Z => n6921);
   U6873 : MUX2_X1 port map( A => REGISTERS_18_2_port, B => n1828, S => n1736, 
                           Z => n6922);
   U6874 : MUX2_X1 port map( A => REGISTERS_18_1_port, B => n1817, S => n1736, 
                           Z => n6923);
   U6875 : MUX2_X1 port map( A => REGISTERS_18_0_port, B => n1806, S => n1736, 
                           Z => n6924);
   U6876 : MUX2_X1 port map( A => REGISTERS_17_31_port, B => n2953, S => n1737,
                           Z => n6861);
   U6877 : MUX2_X1 port map( A => REGISTERS_17_30_port, B => n2942, S => n1737,
                           Z => n6862);
   U6878 : MUX2_X1 port map( A => REGISTERS_17_29_port, B => n2931, S => n1737,
                           Z => n6863);
   U6879 : MUX2_X1 port map( A => REGISTERS_17_28_port, B => n2915, S => n1737,
                           Z => n6864);
   U6880 : MUX2_X1 port map( A => REGISTERS_17_27_port, B => n2904, S => n1737,
                           Z => n6865);
   U6881 : MUX2_X1 port map( A => REGISTERS_17_26_port, B => n2892, S => n1737,
                           Z => n6866);
   U6882 : MUX2_X1 port map( A => REGISTERS_17_25_port, B => n2881, S => n1737,
                           Z => n6867);
   U6883 : MUX2_X1 port map( A => REGISTERS_17_24_port, B => n2870, S => n1737,
                           Z => n6868);
   U6884 : MUX2_X1 port map( A => REGISTERS_17_23_port, B => n2859, S => n1737,
                           Z => n6869);
   U6885 : MUX2_X1 port map( A => REGISTERS_17_22_port, B => n2848, S => n1737,
                           Z => n6870);
   U6886 : MUX2_X1 port map( A => REGISTERS_17_21_port, B => n2837, S => n1737,
                           Z => n6871);
   U6887 : MUX2_X1 port map( A => REGISTERS_17_20_port, B => n2826, S => n1737,
                           Z => n6872);
   U6888 : MUX2_X1 port map( A => REGISTERS_17_19_port, B => n2815, S => n1738,
                           Z => n6873);
   U6889 : MUX2_X1 port map( A => REGISTERS_17_18_port, B => n2804, S => n1738,
                           Z => n6874);
   U6890 : MUX2_X1 port map( A => REGISTERS_17_17_port, B => n2793, S => n1738,
                           Z => n6875);
   U6891 : MUX2_X1 port map( A => REGISTERS_17_16_port, B => n2782, S => n1738,
                           Z => n6876);
   U6892 : MUX2_X1 port map( A => REGISTERS_17_15_port, B => n2771, S => n1738,
                           Z => n6877);
   U6893 : MUX2_X1 port map( A => REGISTERS_17_14_port, B => n2760, S => n1738,
                           Z => n6878);
   U6894 : MUX2_X1 port map( A => REGISTERS_17_13_port, B => n2749, S => n1738,
                           Z => n6879);
   U6895 : MUX2_X1 port map( A => REGISTERS_17_12_port, B => n2738, S => n1738,
                           Z => n6880);
   U6896 : MUX2_X1 port map( A => REGISTERS_17_11_port, B => n2727, S => n1738,
                           Z => n6881);
   U6897 : MUX2_X1 port map( A => REGISTERS_17_10_port, B => n2716, S => n1738,
                           Z => n6882);
   U6898 : MUX2_X1 port map( A => REGISTERS_17_9_port, B => n2705, S => n1738, 
                           Z => n6883);
   U6899 : MUX2_X1 port map( A => REGISTERS_17_8_port, B => n2598, S => n1738, 
                           Z => n6884);
   U6900 : MUX2_X1 port map( A => REGISTERS_17_7_port, B => n2587, S => n1739, 
                           Z => n6885);
   U6901 : MUX2_X1 port map( A => REGISTERS_17_6_port, B => n2576, S => n1739, 
                           Z => n6886);
   U6902 : MUX2_X1 port map( A => REGISTERS_17_5_port, B => n2565, S => n1739, 
                           Z => n6887);
   U6903 : MUX2_X1 port map( A => REGISTERS_17_4_port, B => n2554, S => n1739, 
                           Z => n6888);
   U6904 : MUX2_X1 port map( A => REGISTERS_17_3_port, B => n1839, S => n1739, 
                           Z => n6889);
   U6905 : MUX2_X1 port map( A => REGISTERS_17_2_port, B => n1828, S => n1739, 
                           Z => n6890);
   U6906 : MUX2_X1 port map( A => REGISTERS_17_1_port, B => n1817, S => n1739, 
                           Z => n6891);
   U6907 : MUX2_X1 port map( A => REGISTERS_17_0_port, B => n1806, S => n1739, 
                           Z => n6892);
   U6908 : MUX2_X1 port map( A => REGISTERS_16_31_port, B => n2953, S => n1740,
                           Z => n6829);
   U6909 : MUX2_X1 port map( A => REGISTERS_16_30_port, B => n2942, S => n1740,
                           Z => n6830);
   U6910 : MUX2_X1 port map( A => REGISTERS_16_29_port, B => n2931, S => n1740,
                           Z => n6831);
   U6911 : MUX2_X1 port map( A => REGISTERS_16_28_port, B => n2915, S => n1740,
                           Z => n6832);
   U6912 : MUX2_X1 port map( A => REGISTERS_16_27_port, B => n2904, S => n1740,
                           Z => n6833);
   U6913 : MUX2_X1 port map( A => REGISTERS_16_26_port, B => n2892, S => n1740,
                           Z => n6834);
   U6914 : MUX2_X1 port map( A => REGISTERS_16_25_port, B => n2881, S => n1740,
                           Z => n6835);
   U6915 : MUX2_X1 port map( A => REGISTERS_16_24_port, B => n2870, S => n1740,
                           Z => n6836);
   U6916 : MUX2_X1 port map( A => REGISTERS_16_23_port, B => n2859, S => n1740,
                           Z => n6837);
   U6917 : MUX2_X1 port map( A => REGISTERS_16_22_port, B => n2848, S => n1740,
                           Z => n6838);
   U6918 : MUX2_X1 port map( A => REGISTERS_16_21_port, B => n2837, S => n1740,
                           Z => n6839);
   U6919 : MUX2_X1 port map( A => REGISTERS_16_20_port, B => n2826, S => n1740,
                           Z => n6840);
   U6920 : MUX2_X1 port map( A => REGISTERS_16_19_port, B => n2815, S => n1741,
                           Z => n6841);
   U6921 : MUX2_X1 port map( A => REGISTERS_16_18_port, B => n2804, S => n1741,
                           Z => n6842);
   U6922 : MUX2_X1 port map( A => REGISTERS_16_17_port, B => n2793, S => n1741,
                           Z => n6843);
   U6923 : MUX2_X1 port map( A => REGISTERS_16_16_port, B => n2782, S => n1741,
                           Z => n6844);
   U6924 : MUX2_X1 port map( A => REGISTERS_16_15_port, B => n2771, S => n1741,
                           Z => n6845);
   U6925 : MUX2_X1 port map( A => REGISTERS_16_14_port, B => n2760, S => n1741,
                           Z => n6846);
   U6926 : MUX2_X1 port map( A => REGISTERS_16_13_port, B => n2749, S => n1741,
                           Z => n6847);
   U6927 : MUX2_X1 port map( A => REGISTERS_16_12_port, B => n2738, S => n1741,
                           Z => n6848);
   U6928 : MUX2_X1 port map( A => REGISTERS_16_11_port, B => n2727, S => n1741,
                           Z => n6849);
   U6929 : MUX2_X1 port map( A => REGISTERS_16_10_port, B => n2716, S => n1741,
                           Z => n6850);
   U6930 : MUX2_X1 port map( A => REGISTERS_16_9_port, B => n2705, S => n1741, 
                           Z => n6851);
   U6931 : MUX2_X1 port map( A => REGISTERS_16_8_port, B => n2598, S => n1741, 
                           Z => n6852);
   U6932 : MUX2_X1 port map( A => REGISTERS_16_7_port, B => n2587, S => n1742, 
                           Z => n6853);
   U6933 : MUX2_X1 port map( A => REGISTERS_16_6_port, B => n2576, S => n1742, 
                           Z => n6854);
   U6934 : MUX2_X1 port map( A => REGISTERS_16_5_port, B => n2565, S => n1742, 
                           Z => n6855);
   U6935 : MUX2_X1 port map( A => REGISTERS_16_4_port, B => n2554, S => n1742, 
                           Z => n6856);
   U6936 : MUX2_X1 port map( A => REGISTERS_16_3_port, B => n1839, S => n1742, 
                           Z => n6857);
   U6937 : MUX2_X1 port map( A => REGISTERS_16_2_port, B => n1828, S => n1742, 
                           Z => n6858);
   U6938 : MUX2_X1 port map( A => REGISTERS_16_1_port, B => n1817, S => n1742, 
                           Z => n6859);
   U6939 : MUX2_X1 port map( A => REGISTERS_16_0_port, B => n1806, S => n1742, 
                           Z => n6860);
   U6940 : MUX2_X1 port map( A => n9542, B => n2953, S => n1743, Z => n6797);
   U6941 : MUX2_X1 port map( A => n9543, B => n2942, S => n1743, Z => n6798);
   U6942 : MUX2_X1 port map( A => n9544, B => n2931, S => n1743, Z => n6799);
   U6943 : MUX2_X1 port map( A => n9545, B => n2915, S => n1743, Z => n6800);
   U6944 : MUX2_X1 port map( A => n9546, B => n2904, S => n1743, Z => n6801);
   U6945 : MUX2_X1 port map( A => n9547, B => n2892, S => n1743, Z => n6802);
   U6946 : MUX2_X1 port map( A => n9548, B => n2881, S => n1743, Z => n6803);
   U6947 : MUX2_X1 port map( A => n9549, B => n2870, S => n1743, Z => n6804);
   U6948 : MUX2_X1 port map( A => n9550, B => n2859, S => n1743, Z => n6805);
   U6949 : MUX2_X1 port map( A => n9551, B => n2848, S => n1743, Z => n6806);
   U6950 : MUX2_X1 port map( A => n9552, B => n2837, S => n1743, Z => n6807);
   U6951 : MUX2_X1 port map( A => n9553, B => n2826, S => n1743, Z => n6808);
   U6952 : MUX2_X1 port map( A => n9554, B => n2815, S => n1744, Z => n6809);
   U6953 : MUX2_X1 port map( A => n9555, B => n2804, S => n1744, Z => n6810);
   U6954 : MUX2_X1 port map( A => n9556, B => n2793, S => n1744, Z => n6811);
   U6955 : MUX2_X1 port map( A => n9557, B => n2782, S => n1744, Z => n6812);
   U6956 : MUX2_X1 port map( A => n9558, B => n2771, S => n1744, Z => n6813);
   U6957 : MUX2_X1 port map( A => n9559, B => n2760, S => n1744, Z => n6814);
   U6958 : MUX2_X1 port map( A => n9560, B => n2749, S => n1744, Z => n6815);
   U6959 : MUX2_X1 port map( A => n9561, B => n2738, S => n1744, Z => n6816);
   U6960 : MUX2_X1 port map( A => n9562, B => n2727, S => n1744, Z => n6817);
   U6961 : MUX2_X1 port map( A => n9563, B => n2716, S => n1744, Z => n6818);
   U6962 : MUX2_X1 port map( A => n9564, B => n2705, S => n1744, Z => n6819);
   U6963 : MUX2_X1 port map( A => n9565, B => n2598, S => n1744, Z => n6820);
   U6964 : MUX2_X1 port map( A => n9566, B => n2587, S => n1745, Z => n6821);
   U6965 : MUX2_X1 port map( A => n9567, B => n2576, S => n1745, Z => n6822);
   U6966 : MUX2_X1 port map( A => n9568, B => n2565, S => n1745, Z => n6823);
   U6967 : MUX2_X1 port map( A => n9569, B => n2554, S => n1745, Z => n6824);
   U6968 : MUX2_X1 port map( A => n9570, B => n1839, S => n1745, Z => n6825);
   U6969 : MUX2_X1 port map( A => n9571, B => n1828, S => n1745, Z => n6826);
   U6970 : MUX2_X1 port map( A => n9572, B => n1817, S => n1745, Z => n6827);
   U6971 : MUX2_X1 port map( A => n9573, B => n1806, S => n1745, Z => n6828);
   U6972 : MUX2_X1 port map( A => n9510, B => n2953, S => n1746, Z => n6765);
   U6973 : MUX2_X1 port map( A => n9511, B => n2942, S => n1746, Z => n6766);
   U6974 : MUX2_X1 port map( A => n9512, B => n2931, S => n1746, Z => n6767);
   U6975 : MUX2_X1 port map( A => n9513, B => n2915, S => n1746, Z => n6768);
   U6976 : MUX2_X1 port map( A => n9514, B => n2904, S => n1746, Z => n6769);
   U6977 : MUX2_X1 port map( A => n9515, B => n2892, S => n1746, Z => n6770);
   U6978 : MUX2_X1 port map( A => n9516, B => n2881, S => n1746, Z => n6771);
   U6979 : MUX2_X1 port map( A => n9517, B => n2870, S => n1746, Z => n6772);
   U6980 : MUX2_X1 port map( A => n9518, B => n2859, S => n1746, Z => n6773);
   U6981 : MUX2_X1 port map( A => n9519, B => n2848, S => n1746, Z => n6774);
   U6982 : MUX2_X1 port map( A => n9520, B => n2837, S => n1746, Z => n6775);
   U6983 : MUX2_X1 port map( A => n9521, B => n2826, S => n1746, Z => n6776);
   U6984 : MUX2_X1 port map( A => n9522, B => n2815, S => n1747, Z => n6777);
   U6985 : MUX2_X1 port map( A => n9523, B => n2804, S => n1747, Z => n6778);
   U6986 : MUX2_X1 port map( A => n9524, B => n2793, S => n1747, Z => n6779);
   U6987 : MUX2_X1 port map( A => n9525, B => n2782, S => n1747, Z => n6780);
   U6988 : MUX2_X1 port map( A => n9526, B => n2771, S => n1747, Z => n6781);
   U6989 : MUX2_X1 port map( A => n9527, B => n2760, S => n1747, Z => n6782);
   U6990 : MUX2_X1 port map( A => n9528, B => n2749, S => n1747, Z => n6783);
   U6991 : MUX2_X1 port map( A => n9529, B => n2738, S => n1747, Z => n6784);
   U6992 : MUX2_X1 port map( A => n9530, B => n2727, S => n1747, Z => n6785);
   U6993 : MUX2_X1 port map( A => n9531, B => n2716, S => n1747, Z => n6786);
   U6994 : MUX2_X1 port map( A => n9532, B => n2705, S => n1747, Z => n6787);
   U6995 : MUX2_X1 port map( A => n9533, B => n2598, S => n1747, Z => n6788);
   U6996 : MUX2_X1 port map( A => n9534, B => n2587, S => n1748, Z => n6789);
   U6997 : MUX2_X1 port map( A => n9535, B => n2576, S => n1748, Z => n6790);
   U6998 : MUX2_X1 port map( A => n9536, B => n2565, S => n1748, Z => n6791);
   U6999 : MUX2_X1 port map( A => n9537, B => n2554, S => n1748, Z => n6792);
   U7000 : MUX2_X1 port map( A => n9538, B => n1839, S => n1748, Z => n6793);
   U7001 : MUX2_X1 port map( A => n9539, B => n1828, S => n1748, Z => n6794);
   U7002 : MUX2_X1 port map( A => n9540, B => n1817, S => n1748, Z => n6795);
   U7003 : MUX2_X1 port map( A => n9541, B => n1806, S => n1748, Z => n6796);
   U7004 : MUX2_X1 port map( A => n9478, B => n2953, S => n1749, Z => n6733);
   U7005 : MUX2_X1 port map( A => n9479, B => n2942, S => n1749, Z => n6734);
   U7006 : MUX2_X1 port map( A => n9480, B => n2931, S => n1749, Z => n6735);
   U7007 : MUX2_X1 port map( A => n9481, B => n2915, S => n1749, Z => n6736);
   U7008 : MUX2_X1 port map( A => n9482, B => n2904, S => n1749, Z => n6737);
   U7009 : MUX2_X1 port map( A => n9483, B => n2892, S => n1749, Z => n6738);
   U7010 : MUX2_X1 port map( A => n9484, B => n2881, S => n1749, Z => n6739);
   U7011 : MUX2_X1 port map( A => n9485, B => n2870, S => n1749, Z => n6740);
   U7012 : MUX2_X1 port map( A => n9486, B => n2859, S => n1749, Z => n6741);
   U7013 : MUX2_X1 port map( A => n9487, B => n2848, S => n1749, Z => n6742);
   U7014 : MUX2_X1 port map( A => n9488, B => n2837, S => n1749, Z => n6743);
   U7015 : MUX2_X1 port map( A => n9489, B => n2826, S => n1749, Z => n6744);
   U7016 : MUX2_X1 port map( A => n9490, B => n2815, S => n1750, Z => n6745);
   U7017 : MUX2_X1 port map( A => n9491, B => n2804, S => n1750, Z => n6746);
   U7018 : MUX2_X1 port map( A => n9492, B => n2793, S => n1750, Z => n6747);
   U7019 : MUX2_X1 port map( A => n9493, B => n2782, S => n1750, Z => n6748);
   U7020 : MUX2_X1 port map( A => n9494, B => n2771, S => n1750, Z => n6749);
   U7021 : MUX2_X1 port map( A => n9495, B => n2760, S => n1750, Z => n6750);
   U7022 : MUX2_X1 port map( A => n9496, B => n2749, S => n1750, Z => n6751);
   U7023 : MUX2_X1 port map( A => n9497, B => n2738, S => n1750, Z => n6752);
   U7024 : MUX2_X1 port map( A => n9498, B => n2727, S => n1750, Z => n6753);
   U7025 : MUX2_X1 port map( A => n9499, B => n2716, S => n1750, Z => n6754);
   U7026 : MUX2_X1 port map( A => n9500, B => n2705, S => n1750, Z => n6755);
   U7027 : MUX2_X1 port map( A => n9501, B => n2598, S => n1750, Z => n6756);
   U7028 : MUX2_X1 port map( A => n9502, B => n2587, S => n1751, Z => n6757);
   U7029 : MUX2_X1 port map( A => n9503, B => n2576, S => n1751, Z => n6758);
   U7030 : MUX2_X1 port map( A => n9504, B => n2565, S => n1751, Z => n6759);
   U7031 : MUX2_X1 port map( A => n9505, B => n2554, S => n1751, Z => n6760);
   U7032 : MUX2_X1 port map( A => n9506, B => n1839, S => n1751, Z => n6761);
   U7033 : MUX2_X1 port map( A => n9507, B => n1828, S => n1751, Z => n6762);
   U7034 : MUX2_X1 port map( A => n9508, B => n1817, S => n1751, Z => n6763);
   U7035 : MUX2_X1 port map( A => n9509, B => n1806, S => n1751, Z => n6764);
   U7036 : MUX2_X1 port map( A => REGISTERS_12_31_port, B => n2953, S => n1752,
                           Z => n6701);
   U7037 : MUX2_X1 port map( A => REGISTERS_12_30_port, B => n2942, S => n1752,
                           Z => n6702);
   U7038 : MUX2_X1 port map( A => REGISTERS_12_29_port, B => n2931, S => n1752,
                           Z => n6703);
   U7039 : MUX2_X1 port map( A => REGISTERS_12_28_port, B => n2915, S => n1752,
                           Z => n6704);
   U7040 : MUX2_X1 port map( A => REGISTERS_12_27_port, B => n2904, S => n1752,
                           Z => n6705);
   U7041 : MUX2_X1 port map( A => REGISTERS_12_26_port, B => n2892, S => n1752,
                           Z => n6706);
   U7042 : MUX2_X1 port map( A => REGISTERS_12_25_port, B => n2881, S => n1752,
                           Z => n6707);
   U7043 : MUX2_X1 port map( A => REGISTERS_12_24_port, B => n2870, S => n1752,
                           Z => n6708);
   U7044 : MUX2_X1 port map( A => REGISTERS_12_23_port, B => n2859, S => n1752,
                           Z => n6709);
   U7045 : MUX2_X1 port map( A => REGISTERS_12_22_port, B => n2848, S => n1752,
                           Z => n6710);
   U7046 : MUX2_X1 port map( A => REGISTERS_12_21_port, B => n2837, S => n1752,
                           Z => n6711);
   U7047 : MUX2_X1 port map( A => REGISTERS_12_20_port, B => n2826, S => n1752,
                           Z => n6712);
   U7048 : MUX2_X1 port map( A => REGISTERS_12_19_port, B => n2815, S => n1753,
                           Z => n6713);
   U7049 : MUX2_X1 port map( A => REGISTERS_12_18_port, B => n2804, S => n1753,
                           Z => n6714);
   U7050 : MUX2_X1 port map( A => REGISTERS_12_17_port, B => n2793, S => n1753,
                           Z => n6715);
   U7051 : MUX2_X1 port map( A => REGISTERS_12_16_port, B => n2782, S => n1753,
                           Z => n6716);
   U7052 : MUX2_X1 port map( A => REGISTERS_12_15_port, B => n2771, S => n1753,
                           Z => n6717);
   U7053 : MUX2_X1 port map( A => REGISTERS_12_14_port, B => n2760, S => n1753,
                           Z => n6718);
   U7054 : MUX2_X1 port map( A => REGISTERS_12_13_port, B => n2749, S => n1753,
                           Z => n6719);
   U7055 : MUX2_X1 port map( A => REGISTERS_12_12_port, B => n2738, S => n1753,
                           Z => n6720);
   U7056 : MUX2_X1 port map( A => REGISTERS_12_11_port, B => n2727, S => n1753,
                           Z => n6721);
   U7057 : MUX2_X1 port map( A => REGISTERS_12_10_port, B => n2716, S => n1753,
                           Z => n6722);
   U7058 : MUX2_X1 port map( A => REGISTERS_12_9_port, B => n2705, S => n1753, 
                           Z => n6723);
   U7059 : MUX2_X1 port map( A => REGISTERS_12_8_port, B => n2598, S => n1753, 
                           Z => n6724);
   U7060 : MUX2_X1 port map( A => REGISTERS_12_7_port, B => n2587, S => n1754, 
                           Z => n6725);
   U7061 : MUX2_X1 port map( A => REGISTERS_12_6_port, B => n2576, S => n1754, 
                           Z => n6726);
   U7062 : MUX2_X1 port map( A => REGISTERS_12_5_port, B => n2565, S => n1754, 
                           Z => n6727);
   U7063 : MUX2_X1 port map( A => REGISTERS_12_4_port, B => n2554, S => n1754, 
                           Z => n6728);
   U7064 : MUX2_X1 port map( A => REGISTERS_12_3_port, B => n1839, S => n1754, 
                           Z => n6729);
   U7065 : MUX2_X1 port map( A => REGISTERS_12_2_port, B => n1828, S => n1754, 
                           Z => n6730);
   U7066 : MUX2_X1 port map( A => REGISTERS_12_1_port, B => n1817, S => n1754, 
                           Z => n6731);
   U7067 : MUX2_X1 port map( A => REGISTERS_12_0_port, B => n1806, S => n1754, 
                           Z => n6732);
   U7068 : MUX2_X1 port map( A => REGISTERS_11_31_port, B => n2953, S => n1755,
                           Z => n6669);
   U7069 : MUX2_X1 port map( A => REGISTERS_11_30_port, B => n2942, S => n1755,
                           Z => n6670);
   U7070 : MUX2_X1 port map( A => REGISTERS_11_29_port, B => n2931, S => n1755,
                           Z => n6671);
   U7071 : MUX2_X1 port map( A => REGISTERS_11_28_port, B => n2915, S => n1755,
                           Z => n6672);
   U7072 : MUX2_X1 port map( A => REGISTERS_11_27_port, B => n2904, S => n1755,
                           Z => n6673);
   U7073 : MUX2_X1 port map( A => REGISTERS_11_26_port, B => n2892, S => n1755,
                           Z => n6674);
   U7074 : MUX2_X1 port map( A => REGISTERS_11_25_port, B => n2881, S => n1755,
                           Z => n6675);
   U7075 : MUX2_X1 port map( A => REGISTERS_11_24_port, B => n2870, S => n1755,
                           Z => n6676);
   U7076 : MUX2_X1 port map( A => REGISTERS_11_23_port, B => n2859, S => n1755,
                           Z => n6677);
   U7077 : MUX2_X1 port map( A => REGISTERS_11_22_port, B => n2848, S => n1755,
                           Z => n6678);
   U7078 : MUX2_X1 port map( A => REGISTERS_11_21_port, B => n2837, S => n1755,
                           Z => n6679);
   U7079 : MUX2_X1 port map( A => REGISTERS_11_20_port, B => n2826, S => n1755,
                           Z => n6680);
   U7080 : MUX2_X1 port map( A => REGISTERS_11_19_port, B => n2815, S => n1756,
                           Z => n6681);
   U7081 : MUX2_X1 port map( A => REGISTERS_11_18_port, B => n2804, S => n1756,
                           Z => n6682);
   U7082 : MUX2_X1 port map( A => REGISTERS_11_17_port, B => n2793, S => n1756,
                           Z => n6683);
   U7083 : MUX2_X1 port map( A => REGISTERS_11_16_port, B => n2782, S => n1756,
                           Z => n6684);
   U7084 : MUX2_X1 port map( A => REGISTERS_11_15_port, B => n2771, S => n1756,
                           Z => n6685);
   U7085 : MUX2_X1 port map( A => REGISTERS_11_14_port, B => n2760, S => n1756,
                           Z => n6686);
   U7086 : MUX2_X1 port map( A => REGISTERS_11_13_port, B => n2749, S => n1756,
                           Z => n6687);
   U7087 : MUX2_X1 port map( A => REGISTERS_11_12_port, B => n2738, S => n1756,
                           Z => n6688);
   U7088 : MUX2_X1 port map( A => REGISTERS_11_11_port, B => n2727, S => n1756,
                           Z => n6689);
   U7089 : MUX2_X1 port map( A => REGISTERS_11_10_port, B => n2716, S => n1756,
                           Z => n6690);
   U7090 : MUX2_X1 port map( A => REGISTERS_11_9_port, B => n2705, S => n1756, 
                           Z => n6691);
   U7091 : MUX2_X1 port map( A => REGISTERS_11_8_port, B => n2598, S => n1756, 
                           Z => n6692);
   U7092 : MUX2_X1 port map( A => REGISTERS_11_7_port, B => n2587, S => n1757, 
                           Z => n6693);
   U7093 : MUX2_X1 port map( A => REGISTERS_11_6_port, B => n2576, S => n1757, 
                           Z => n6694);
   U7094 : MUX2_X1 port map( A => REGISTERS_11_5_port, B => n2565, S => n1757, 
                           Z => n6695);
   U7095 : MUX2_X1 port map( A => REGISTERS_11_4_port, B => n2554, S => n1757, 
                           Z => n6696);
   U7096 : MUX2_X1 port map( A => REGISTERS_11_3_port, B => n1839, S => n1757, 
                           Z => n6697);
   U7097 : MUX2_X1 port map( A => REGISTERS_11_2_port, B => n1828, S => n1757, 
                           Z => n6698);
   U7098 : MUX2_X1 port map( A => REGISTERS_11_1_port, B => n1817, S => n1757, 
                           Z => n6699);
   U7099 : MUX2_X1 port map( A => REGISTERS_11_0_port, B => n1806, S => n1757, 
                           Z => n6700);
   U7100 : MUX2_X1 port map( A => n9446, B => n2954, S => n1758, Z => n6637);
   U7101 : MUX2_X1 port map( A => n9447, B => n2943, S => n1758, Z => n6638);
   U7102 : MUX2_X1 port map( A => n9448, B => n2932, S => n1758, Z => n6639);
   U7103 : MUX2_X1 port map( A => n9449, B => n2917, S => n1758, Z => n6640);
   U7104 : MUX2_X1 port map( A => n9450, B => n2905, S => n1758, Z => n6641);
   U7105 : MUX2_X1 port map( A => n9451, B => n2893, S => n1758, Z => n6642);
   U7106 : MUX2_X1 port map( A => n9452, B => n2882, S => n1758, Z => n6643);
   U7107 : MUX2_X1 port map( A => n9453, B => n2871, S => n1758, Z => n6644);
   U7108 : MUX2_X1 port map( A => n9454, B => n2860, S => n1758, Z => n6645);
   U7109 : MUX2_X1 port map( A => n9455, B => n2849, S => n1758, Z => n6646);
   U7110 : MUX2_X1 port map( A => n9456, B => n2838, S => n1758, Z => n6647);
   U7111 : MUX2_X1 port map( A => n9457, B => n2827, S => n1758, Z => n6648);
   U7112 : MUX2_X1 port map( A => n9458, B => n2816, S => n1759, Z => n6649);
   U7113 : MUX2_X1 port map( A => n9459, B => n2805, S => n1759, Z => n6650);
   U7114 : MUX2_X1 port map( A => n9460, B => n2794, S => n1759, Z => n6651);
   U7115 : MUX2_X1 port map( A => n9461, B => n2783, S => n1759, Z => n6652);
   U7116 : MUX2_X1 port map( A => n9462, B => n2772, S => n1759, Z => n6653);
   U7117 : MUX2_X1 port map( A => n9463, B => n2761, S => n1759, Z => n6654);
   U7118 : MUX2_X1 port map( A => n9464, B => n2750, S => n1759, Z => n6655);
   U7119 : MUX2_X1 port map( A => n9465, B => n2739, S => n1759, Z => n6656);
   U7120 : MUX2_X1 port map( A => n9466, B => n2728, S => n1759, Z => n6657);
   U7121 : MUX2_X1 port map( A => n9467, B => n2717, S => n1759, Z => n6658);
   U7122 : MUX2_X1 port map( A => n9468, B => n2706, S => n1759, Z => n6659);
   U7123 : MUX2_X1 port map( A => n9469, B => n2599, S => n1759, Z => n6660);
   U7124 : MUX2_X1 port map( A => n9470, B => n2588, S => n1760, Z => n6661);
   U7125 : MUX2_X1 port map( A => n9471, B => n2577, S => n1760, Z => n6662);
   U7126 : MUX2_X1 port map( A => n9472, B => n2566, S => n1760, Z => n6663);
   U7127 : MUX2_X1 port map( A => n9473, B => n2555, S => n1760, Z => n6664);
   U7128 : MUX2_X1 port map( A => n9474, B => n2544, S => n1760, Z => n6665);
   U7129 : MUX2_X1 port map( A => n9475, B => n1829, S => n1760, Z => n6666);
   U7130 : MUX2_X1 port map( A => n9476, B => n1818, S => n1760, Z => n6667);
   U7131 : MUX2_X1 port map( A => n9477, B => n1807, S => n1760, Z => n6668);
   U7132 : MUX2_X1 port map( A => n9414, B => n2954, S => n1761, Z => n6605);
   U7133 : MUX2_X1 port map( A => n9415, B => n2943, S => n1761, Z => n6606);
   U7134 : MUX2_X1 port map( A => n9416, B => n2932, S => n1761, Z => n6607);
   U7135 : MUX2_X1 port map( A => n9417, B => n2917, S => n1761, Z => n6608);
   U7136 : MUX2_X1 port map( A => n9418, B => n2905, S => n1761, Z => n6609);
   U7137 : MUX2_X1 port map( A => n9419, B => n2893, S => n1761, Z => n6610);
   U7138 : MUX2_X1 port map( A => n9420, B => n2882, S => n1761, Z => n6611);
   U7139 : MUX2_X1 port map( A => n9421, B => n2871, S => n1761, Z => n6612);
   U7140 : MUX2_X1 port map( A => n9422, B => n2860, S => n1761, Z => n6613);
   U7141 : MUX2_X1 port map( A => n9423, B => n2849, S => n1761, Z => n6614);
   U7142 : MUX2_X1 port map( A => n9424, B => n2838, S => n1761, Z => n6615);
   U7143 : MUX2_X1 port map( A => n9425, B => n2827, S => n1761, Z => n6616);
   U7144 : MUX2_X1 port map( A => n9426, B => n2816, S => n1762, Z => n6617);
   U7145 : MUX2_X1 port map( A => n9427, B => n2805, S => n1762, Z => n6618);
   U7146 : MUX2_X1 port map( A => n9428, B => n2794, S => n1762, Z => n6619);
   U7147 : MUX2_X1 port map( A => n9429, B => n2783, S => n1762, Z => n6620);
   U7148 : MUX2_X1 port map( A => n9430, B => n2772, S => n1762, Z => n6621);
   U7149 : MUX2_X1 port map( A => n9431, B => n2761, S => n1762, Z => n6622);
   U7150 : MUX2_X1 port map( A => n9432, B => n2750, S => n1762, Z => n6623);
   U7151 : MUX2_X1 port map( A => n9433, B => n2739, S => n1762, Z => n6624);
   U7152 : MUX2_X1 port map( A => n9434, B => n2728, S => n1762, Z => n6625);
   U7153 : MUX2_X1 port map( A => n9435, B => n2717, S => n1762, Z => n6626);
   U7154 : MUX2_X1 port map( A => n9436, B => n2706, S => n1762, Z => n6627);
   U7155 : MUX2_X1 port map( A => n9437, B => n2599, S => n1762, Z => n6628);
   U7156 : MUX2_X1 port map( A => n9438, B => n2588, S => n1763, Z => n6629);
   U7157 : MUX2_X1 port map( A => n9439, B => n2577, S => n1763, Z => n6630);
   U7158 : MUX2_X1 port map( A => n9440, B => n2566, S => n1763, Z => n6631);
   U7159 : MUX2_X1 port map( A => n9441, B => n2555, S => n1763, Z => n6632);
   U7160 : MUX2_X1 port map( A => n9442, B => n2544, S => n1763, Z => n6633);
   U7161 : MUX2_X1 port map( A => n9443, B => n1829, S => n1763, Z => n6634);
   U7162 : MUX2_X1 port map( A => n9444, B => n1818, S => n1763, Z => n6635);
   U7163 : MUX2_X1 port map( A => n9445, B => n1807, S => n1763, Z => n6636);
   U7164 : MUX2_X1 port map( A => n9382, B => n2954, S => n1764, Z => n6573);
   U7165 : MUX2_X1 port map( A => n9383, B => n2943, S => n1764, Z => n6574);
   U7166 : MUX2_X1 port map( A => n9384, B => n2932, S => n1764, Z => n6575);
   U7167 : MUX2_X1 port map( A => n9385, B => n2917, S => n1764, Z => n6576);
   U7168 : MUX2_X1 port map( A => n9386, B => n2905, S => n1764, Z => n6577);
   U7169 : MUX2_X1 port map( A => n9387, B => n2893, S => n1764, Z => n6578);
   U7170 : MUX2_X1 port map( A => n9388, B => n2882, S => n1764, Z => n6579);
   U7171 : MUX2_X1 port map( A => n9389, B => n2871, S => n1764, Z => n6580);
   U7172 : MUX2_X1 port map( A => n9390, B => n2860, S => n1764, Z => n6581);
   U7173 : MUX2_X1 port map( A => n9391, B => n2849, S => n1764, Z => n6582);
   U7174 : MUX2_X1 port map( A => n9392, B => n2838, S => n1764, Z => n6583);
   U7175 : MUX2_X1 port map( A => n9393, B => n2827, S => n1764, Z => n6584);
   U7176 : MUX2_X1 port map( A => n9394, B => n2816, S => n1765, Z => n6585);
   U7177 : MUX2_X1 port map( A => n9395, B => n2805, S => n1765, Z => n6586);
   U7178 : MUX2_X1 port map( A => n9396, B => n2794, S => n1765, Z => n6587);
   U7179 : MUX2_X1 port map( A => n9397, B => n2783, S => n1765, Z => n6588);
   U7180 : MUX2_X1 port map( A => n9398, B => n2772, S => n1765, Z => n6589);
   U7181 : MUX2_X1 port map( A => n9399, B => n2761, S => n1765, Z => n6590);
   U7182 : MUX2_X1 port map( A => n9400, B => n2750, S => n1765, Z => n6591);
   U7183 : MUX2_X1 port map( A => n9401, B => n2739, S => n1765, Z => n6592);
   U7184 : MUX2_X1 port map( A => n9402, B => n2728, S => n1765, Z => n6593);
   U7185 : MUX2_X1 port map( A => n9403, B => n2717, S => n1765, Z => n6594);
   U7186 : MUX2_X1 port map( A => n9404, B => n2706, S => n1765, Z => n6595);
   U7187 : MUX2_X1 port map( A => n9405, B => n2599, S => n1765, Z => n6596);
   U7188 : MUX2_X1 port map( A => n9406, B => n2588, S => n1766, Z => n6597);
   U7189 : MUX2_X1 port map( A => n9407, B => n2577, S => n1766, Z => n6598);
   U7190 : MUX2_X1 port map( A => n9408, B => n2566, S => n1766, Z => n6599);
   U7191 : MUX2_X1 port map( A => n9409, B => n2555, S => n1766, Z => n6600);
   U7192 : MUX2_X1 port map( A => n9410, B => n2544, S => n1766, Z => n6601);
   U7193 : MUX2_X1 port map( A => n9411, B => n1829, S => n1766, Z => n6602);
   U7194 : MUX2_X1 port map( A => n9412, B => n1818, S => n1766, Z => n6603);
   U7195 : MUX2_X1 port map( A => n9413, B => n1807, S => n1766, Z => n6604);
   U7196 : MUX2_X1 port map( A => n9350, B => n2954, S => n1767, Z => n6541);
   U7197 : MUX2_X1 port map( A => n9351, B => n2943, S => n1767, Z => n6542);
   U7198 : MUX2_X1 port map( A => n9352, B => n2932, S => n1767, Z => n6543);
   U7199 : MUX2_X1 port map( A => n9353, B => n2917, S => n1767, Z => n6544);
   U7200 : MUX2_X1 port map( A => n9354, B => n2905, S => n1767, Z => n6545);
   U7201 : MUX2_X1 port map( A => n9355, B => n2893, S => n1767, Z => n6546);
   U7202 : MUX2_X1 port map( A => n9356, B => n2882, S => n1767, Z => n6547);
   U7203 : MUX2_X1 port map( A => n9357, B => n2871, S => n1767, Z => n6548);
   U7204 : MUX2_X1 port map( A => n9358, B => n2860, S => n1767, Z => n6549);
   U7205 : MUX2_X1 port map( A => n9359, B => n2849, S => n1767, Z => n6550);
   U7206 : MUX2_X1 port map( A => n9360, B => n2838, S => n1767, Z => n6551);
   U7207 : MUX2_X1 port map( A => n9361, B => n2827, S => n1767, Z => n6552);
   U7208 : MUX2_X1 port map( A => n9362, B => n2816, S => n1768, Z => n6553);
   U7209 : MUX2_X1 port map( A => n9363, B => n2805, S => n1768, Z => n6554);
   U7210 : MUX2_X1 port map( A => n9364, B => n2794, S => n1768, Z => n6555);
   U7211 : MUX2_X1 port map( A => n9365, B => n2783, S => n1768, Z => n6556);
   U7212 : MUX2_X1 port map( A => n9366, B => n2772, S => n1768, Z => n6557);
   U7213 : MUX2_X1 port map( A => n9367, B => n2761, S => n1768, Z => n6558);
   U7214 : MUX2_X1 port map( A => n9368, B => n2750, S => n1768, Z => n6559);
   U7215 : MUX2_X1 port map( A => n9369, B => n2739, S => n1768, Z => n6560);
   U7216 : MUX2_X1 port map( A => n9370, B => n2728, S => n1768, Z => n6561);
   U7217 : MUX2_X1 port map( A => n9371, B => n2717, S => n1768, Z => n6562);
   U7218 : MUX2_X1 port map( A => n9372, B => n2706, S => n1768, Z => n6563);
   U7219 : MUX2_X1 port map( A => n9373, B => n2599, S => n1768, Z => n6564);
   U7220 : MUX2_X1 port map( A => n9374, B => n2588, S => n1769, Z => n6565);
   U7221 : MUX2_X1 port map( A => n9375, B => n2577, S => n1769, Z => n6566);
   U7222 : MUX2_X1 port map( A => n9376, B => n2566, S => n1769, Z => n6567);
   U7223 : MUX2_X1 port map( A => n9377, B => n2555, S => n1769, Z => n6568);
   U7224 : MUX2_X1 port map( A => n9378, B => n2544, S => n1769, Z => n6569);
   U7225 : MUX2_X1 port map( A => n9379, B => n1829, S => n1769, Z => n6570);
   U7226 : MUX2_X1 port map( A => n9380, B => n1818, S => n1769, Z => n6571);
   U7227 : MUX2_X1 port map( A => n9381, B => n1807, S => n1769, Z => n6572);
   U7228 : MUX2_X1 port map( A => n9318, B => n2954, S => n1770, Z => n6509);
   U7229 : MUX2_X1 port map( A => n9319, B => n2943, S => n1770, Z => n6510);
   U7230 : MUX2_X1 port map( A => n9320, B => n2932, S => n1770, Z => n6511);
   U7231 : MUX2_X1 port map( A => n9321, B => n2917, S => n1770, Z => n6512);
   U7232 : MUX2_X1 port map( A => n9322, B => n2905, S => n1770, Z => n6513);
   U7233 : MUX2_X1 port map( A => n9323, B => n2893, S => n1770, Z => n6514);
   U7234 : MUX2_X1 port map( A => n9324, B => n2882, S => n1770, Z => n6515);
   U7235 : MUX2_X1 port map( A => n9325, B => n2871, S => n1770, Z => n6516);
   U7236 : MUX2_X1 port map( A => n9326, B => n2860, S => n1770, Z => n6517);
   U7237 : MUX2_X1 port map( A => n9327, B => n2849, S => n1770, Z => n6518);
   U7238 : MUX2_X1 port map( A => n9328, B => n2838, S => n1770, Z => n6519);
   U7239 : MUX2_X1 port map( A => n9329, B => n2827, S => n1770, Z => n6520);
   U7240 : MUX2_X1 port map( A => n9330, B => n2816, S => n1771, Z => n6521);
   U7241 : MUX2_X1 port map( A => n9331, B => n2805, S => n1771, Z => n6522);
   U7242 : MUX2_X1 port map( A => n9332, B => n2794, S => n1771, Z => n6523);
   U7243 : MUX2_X1 port map( A => n9333, B => n2783, S => n1771, Z => n6524);
   U7244 : MUX2_X1 port map( A => n9334, B => n2772, S => n1771, Z => n6525);
   U7245 : MUX2_X1 port map( A => n9335, B => n2761, S => n1771, Z => n6526);
   U7246 : MUX2_X1 port map( A => n9336, B => n2750, S => n1771, Z => n6527);
   U7247 : MUX2_X1 port map( A => n9337, B => n2739, S => n1771, Z => n6528);
   U7248 : MUX2_X1 port map( A => n9338, B => n2728, S => n1771, Z => n6529);
   U7249 : MUX2_X1 port map( A => n9339, B => n2717, S => n1771, Z => n6530);
   U7250 : MUX2_X1 port map( A => n9340, B => n2706, S => n1771, Z => n6531);
   U7251 : MUX2_X1 port map( A => n9341, B => n2599, S => n1771, Z => n6532);
   U7252 : MUX2_X1 port map( A => n9342, B => n2588, S => n1772, Z => n6533);
   U7253 : MUX2_X1 port map( A => n9343, B => n2577, S => n1772, Z => n6534);
   U7254 : MUX2_X1 port map( A => n9344, B => n2566, S => n1772, Z => n6535);
   U7255 : MUX2_X1 port map( A => n9345, B => n2555, S => n1772, Z => n6536);
   U7256 : MUX2_X1 port map( A => n9346, B => n2544, S => n1772, Z => n6537);
   U7257 : MUX2_X1 port map( A => n9347, B => n1829, S => n1772, Z => n6538);
   U7258 : MUX2_X1 port map( A => n9348, B => n1818, S => n1772, Z => n6539);
   U7259 : MUX2_X1 port map( A => n9349, B => n1807, S => n1772, Z => n6540);
   U7260 : MUX2_X1 port map( A => n9286, B => n2954, S => n1773, Z => n6477);
   U7261 : MUX2_X1 port map( A => n9287, B => n2943, S => n1773, Z => n6478);
   U7262 : MUX2_X1 port map( A => n9288, B => n2932, S => n1773, Z => n6479);
   U7263 : MUX2_X1 port map( A => n9289, B => n2917, S => n1773, Z => n6480);
   U7264 : MUX2_X1 port map( A => n9290, B => n2905, S => n1773, Z => n6481);
   U7265 : MUX2_X1 port map( A => n9291, B => n2893, S => n1773, Z => n6482);
   U7266 : MUX2_X1 port map( A => n9292, B => n2882, S => n1773, Z => n6483);
   U7267 : MUX2_X1 port map( A => n9293, B => n2871, S => n1773, Z => n6484);
   U7268 : MUX2_X1 port map( A => n9294, B => n2860, S => n1773, Z => n6485);
   U7269 : MUX2_X1 port map( A => n9295, B => n2849, S => n1773, Z => n6486);
   U7270 : MUX2_X1 port map( A => n9296, B => n2838, S => n1773, Z => n6487);
   U7271 : MUX2_X1 port map( A => n9297, B => n2827, S => n1773, Z => n6488);
   U7272 : MUX2_X1 port map( A => n9298, B => n2816, S => n1774, Z => n6489);
   U7273 : MUX2_X1 port map( A => n9299, B => n2805, S => n1774, Z => n6490);
   U7274 : MUX2_X1 port map( A => n9300, B => n2794, S => n1774, Z => n6491);
   U7275 : MUX2_X1 port map( A => n9301, B => n2783, S => n1774, Z => n6492);
   U7276 : MUX2_X1 port map( A => n9302, B => n2772, S => n1774, Z => n6493);
   U7277 : MUX2_X1 port map( A => n9303, B => n2761, S => n1774, Z => n6494);
   U7278 : MUX2_X1 port map( A => n9304, B => n2750, S => n1774, Z => n6495);
   U7279 : MUX2_X1 port map( A => n9305, B => n2739, S => n1774, Z => n6496);
   U7280 : MUX2_X1 port map( A => n9306, B => n2728, S => n1774, Z => n6497);
   U7281 : MUX2_X1 port map( A => n9307, B => n2717, S => n1774, Z => n6498);
   U7282 : MUX2_X1 port map( A => n9308, B => n2706, S => n1774, Z => n6499);
   U7283 : MUX2_X1 port map( A => n9309, B => n2599, S => n1774, Z => n6500);
   U7284 : MUX2_X1 port map( A => n9310, B => n2588, S => n1775, Z => n6501);
   U7285 : MUX2_X1 port map( A => n9311, B => n2577, S => n1775, Z => n6502);
   U7286 : MUX2_X1 port map( A => n9312, B => n2566, S => n1775, Z => n6503);
   U7287 : MUX2_X1 port map( A => n9313, B => n2555, S => n1775, Z => n6504);
   U7288 : MUX2_X1 port map( A => n9314, B => n2544, S => n1775, Z => n6505);
   U7289 : MUX2_X1 port map( A => n9315, B => n1829, S => n1775, Z => n6506);
   U7290 : MUX2_X1 port map( A => n9316, B => n1818, S => n1775, Z => n6507);
   U7291 : MUX2_X1 port map( A => n9317, B => n1807, S => n1775, Z => n6508);
   U7292 : MUX2_X1 port map( A => n9254, B => n2954, S => n1776, Z => n6445);
   U7293 : MUX2_X1 port map( A => n9255, B => n2943, S => n1776, Z => n6446);
   U7294 : MUX2_X1 port map( A => n9256, B => n2932, S => n1776, Z => n6447);
   U7295 : MUX2_X1 port map( A => n9257, B => n2917, S => n1776, Z => n6448);
   U7296 : MUX2_X1 port map( A => n9258, B => n2905, S => n1776, Z => n6449);
   U7297 : MUX2_X1 port map( A => n9259, B => n2893, S => n1776, Z => n6450);
   U7298 : MUX2_X1 port map( A => n9260, B => n2882, S => n1776, Z => n6451);
   U7299 : MUX2_X1 port map( A => n9261, B => n2871, S => n1776, Z => n6452);
   U7300 : MUX2_X1 port map( A => n9262, B => n2860, S => n1776, Z => n6453);
   U7301 : MUX2_X1 port map( A => n9263, B => n2849, S => n1776, Z => n6454);
   U7302 : MUX2_X1 port map( A => n9264, B => n2838, S => n1776, Z => n6455);
   U7303 : MUX2_X1 port map( A => n9265, B => n2827, S => n1776, Z => n6456);
   U7304 : MUX2_X1 port map( A => n9266, B => n2816, S => n1777, Z => n6457);
   U7305 : MUX2_X1 port map( A => n9267, B => n2805, S => n1777, Z => n6458);
   U7306 : MUX2_X1 port map( A => n9268, B => n2794, S => n1777, Z => n6459);
   U7307 : MUX2_X1 port map( A => n9269, B => n2783, S => n1777, Z => n6460);
   U7308 : MUX2_X1 port map( A => n9270, B => n2772, S => n1777, Z => n6461);
   U7309 : MUX2_X1 port map( A => n9271, B => n2761, S => n1777, Z => n6462);
   U7310 : MUX2_X1 port map( A => n9272, B => n2750, S => n1777, Z => n6463);
   U7311 : MUX2_X1 port map( A => n9273, B => n2739, S => n1777, Z => n6464);
   U7312 : MUX2_X1 port map( A => n9274, B => n2728, S => n1777, Z => n6465);
   U7313 : MUX2_X1 port map( A => n9275, B => n2717, S => n1777, Z => n6466);
   U7314 : MUX2_X1 port map( A => n9276, B => n2706, S => n1777, Z => n6467);
   U7315 : MUX2_X1 port map( A => n9277, B => n2599, S => n1777, Z => n6468);
   U7316 : MUX2_X1 port map( A => n9278, B => n2588, S => n1778, Z => n6469);
   U7317 : MUX2_X1 port map( A => n9279, B => n2577, S => n1778, Z => n6470);
   U7318 : MUX2_X1 port map( A => n9280, B => n2566, S => n1778, Z => n6471);
   U7319 : MUX2_X1 port map( A => n9281, B => n2555, S => n1778, Z => n6472);
   U7320 : MUX2_X1 port map( A => n9282, B => n2544, S => n1778, Z => n6473);
   U7321 : MUX2_X1 port map( A => n9283, B => n1829, S => n1778, Z => n6474);
   U7322 : MUX2_X1 port map( A => n9284, B => n1818, S => n1778, Z => n6475);
   U7323 : MUX2_X1 port map( A => n9285, B => n1807, S => n1778, Z => n6476);
   U7324 : MUX2_X1 port map( A => n9222, B => n2954, S => n1779, Z => n6413);
   U7325 : MUX2_X1 port map( A => n9223, B => n2943, S => n1779, Z => n6414);
   U7326 : MUX2_X1 port map( A => n9224, B => n2932, S => n1779, Z => n6415);
   U7327 : MUX2_X1 port map( A => n9225, B => n2917, S => n1779, Z => n6416);
   U7328 : MUX2_X1 port map( A => n9226, B => n2905, S => n1779, Z => n6417);
   U7329 : MUX2_X1 port map( A => n9227, B => n2893, S => n1779, Z => n6418);
   U7330 : MUX2_X1 port map( A => n9228, B => n2882, S => n1779, Z => n6419);
   U7331 : MUX2_X1 port map( A => n9229, B => n2871, S => n1779, Z => n6420);
   U7332 : MUX2_X1 port map( A => n9230, B => n2860, S => n1779, Z => n6421);
   U7333 : MUX2_X1 port map( A => n9231, B => n2849, S => n1779, Z => n6422);
   U7334 : MUX2_X1 port map( A => n9232, B => n2838, S => n1779, Z => n6423);
   U7335 : MUX2_X1 port map( A => n9233, B => n2827, S => n1779, Z => n6424);
   U7336 : MUX2_X1 port map( A => n9234, B => n2816, S => n1780, Z => n6425);
   U7337 : MUX2_X1 port map( A => n9235, B => n2805, S => n1780, Z => n6426);
   U7338 : MUX2_X1 port map( A => n9236, B => n2794, S => n1780, Z => n6427);
   U7339 : MUX2_X1 port map( A => n9237, B => n2783, S => n1780, Z => n6428);
   U7340 : MUX2_X1 port map( A => n9238, B => n2772, S => n1780, Z => n6429);
   U7341 : MUX2_X1 port map( A => n9239, B => n2761, S => n1780, Z => n6430);
   U7342 : MUX2_X1 port map( A => n9240, B => n2750, S => n1780, Z => n6431);
   U7343 : MUX2_X1 port map( A => n9241, B => n2739, S => n1780, Z => n6432);
   U7344 : MUX2_X1 port map( A => n9242, B => n2728, S => n1780, Z => n6433);
   U7345 : MUX2_X1 port map( A => n9243, B => n2717, S => n1780, Z => n6434);
   U7346 : MUX2_X1 port map( A => n9244, B => n2706, S => n1780, Z => n6435);
   U7347 : MUX2_X1 port map( A => n9245, B => n2599, S => n1780, Z => n6436);
   U7348 : MUX2_X1 port map( A => n9246, B => n2588, S => n1781, Z => n6437);
   U7349 : MUX2_X1 port map( A => n9247, B => n2577, S => n1781, Z => n6438);
   U7350 : MUX2_X1 port map( A => n9248, B => n2566, S => n1781, Z => n6439);
   U7351 : MUX2_X1 port map( A => n9249, B => n2555, S => n1781, Z => n6440);
   U7352 : MUX2_X1 port map( A => n9250, B => n2544, S => n1781, Z => n6441);
   U7353 : MUX2_X1 port map( A => n9251, B => n1829, S => n1781, Z => n6442);
   U7354 : MUX2_X1 port map( A => n9252, B => n1818, S => n1781, Z => n6443);
   U7355 : MUX2_X1 port map( A => n9253, B => n1807, S => n1781, Z => n6444);
   U7356 : MUX2_X1 port map( A => n9190, B => n2954, S => n1782, Z => n6381);
   U7357 : MUX2_X1 port map( A => n9191, B => n2943, S => n1782, Z => n6382);
   U7358 : MUX2_X1 port map( A => n9192, B => n2932, S => n1782, Z => n6383);
   U7359 : MUX2_X1 port map( A => n9193, B => n2917, S => n1782, Z => n6384);
   U7360 : MUX2_X1 port map( A => n9194, B => n2905, S => n1782, Z => n6385);
   U7361 : MUX2_X1 port map( A => n9195, B => n2893, S => n1782, Z => n6386);
   U7362 : MUX2_X1 port map( A => n9196, B => n2882, S => n1782, Z => n6387);
   U7363 : MUX2_X1 port map( A => n9197, B => n2871, S => n1782, Z => n6388);
   U7364 : MUX2_X1 port map( A => n9198, B => n2860, S => n1782, Z => n6389);
   U7365 : MUX2_X1 port map( A => n9199, B => n2849, S => n1782, Z => n6390);
   U7366 : MUX2_X1 port map( A => n9200, B => n2838, S => n1782, Z => n6391);
   U7367 : MUX2_X1 port map( A => n9201, B => n2827, S => n1782, Z => n6392);
   U7368 : MUX2_X1 port map( A => n9202, B => n2816, S => n1783, Z => n6393);
   U7369 : MUX2_X1 port map( A => n9203, B => n2805, S => n1783, Z => n6394);
   U7370 : MUX2_X1 port map( A => n9204, B => n2794, S => n1783, Z => n6395);
   U7371 : MUX2_X1 port map( A => n9205, B => n2783, S => n1783, Z => n6396);
   U7372 : MUX2_X1 port map( A => n9206, B => n2772, S => n1783, Z => n6397);
   U7373 : MUX2_X1 port map( A => n9207, B => n2761, S => n1783, Z => n6398);
   U7374 : MUX2_X1 port map( A => n9208, B => n2750, S => n1783, Z => n6399);
   U7375 : MUX2_X1 port map( A => n9209, B => n2739, S => n1783, Z => n6400);
   U7376 : MUX2_X1 port map( A => n9210, B => n2728, S => n1783, Z => n6401);
   U7377 : MUX2_X1 port map( A => n9211, B => n2717, S => n1783, Z => n6402);
   U7378 : MUX2_X1 port map( A => n9212, B => n2706, S => n1783, Z => n6403);
   U7379 : MUX2_X1 port map( A => n9213, B => n2599, S => n1783, Z => n6404);
   U7380 : MUX2_X1 port map( A => n9214, B => n2588, S => n1784, Z => n6405);
   U7381 : MUX2_X1 port map( A => n9215, B => n2577, S => n1784, Z => n6406);
   U7382 : MUX2_X1 port map( A => n9216, B => n2566, S => n1784, Z => n6407);
   U7383 : MUX2_X1 port map( A => n9217, B => n2555, S => n1784, Z => n6408);
   U7384 : MUX2_X1 port map( A => n9218, B => n2544, S => n1784, Z => n6409);
   U7385 : MUX2_X1 port map( A => n9219, B => n1829, S => n1784, Z => n6410);
   U7386 : MUX2_X1 port map( A => n9220, B => n1818, S => n1784, Z => n6411);
   U7387 : MUX2_X1 port map( A => n9221, B => n1807, S => n1784, Z => n6412);
   U7388 : MUX2_X1 port map( A => n9158, B => n2954, S => n1785, Z => n6349);
   U7389 : MUX2_X1 port map( A => n9159, B => n2943, S => n1785, Z => n6350);
   U7390 : MUX2_X1 port map( A => n9160, B => n2932, S => n1785, Z => n6351);
   U7391 : MUX2_X1 port map( A => n9161, B => n2917, S => n1785, Z => n6352);
   U7392 : MUX2_X1 port map( A => n9162, B => n2905, S => n1785, Z => n6353);
   U7393 : MUX2_X1 port map( A => n9163, B => n2893, S => n1785, Z => n6354);
   U7394 : MUX2_X1 port map( A => n9164, B => n2882, S => n1785, Z => n6355);
   U7395 : MUX2_X1 port map( A => n9165, B => n2871, S => n1785, Z => n6356);
   U7396 : MUX2_X1 port map( A => n9166, B => n2860, S => n1785, Z => n6357);
   U7397 : MUX2_X1 port map( A => n9167, B => n2849, S => n1785, Z => n6358);
   U7398 : MUX2_X1 port map( A => n9168, B => n2838, S => n1785, Z => n6359);
   U7399 : MUX2_X1 port map( A => n9169, B => n2827, S => n1785, Z => n6360);
   U7400 : MUX2_X1 port map( A => n9170, B => n2816, S => n1786, Z => n6361);
   U7401 : MUX2_X1 port map( A => n9171, B => n2805, S => n1786, Z => n6362);
   U7402 : MUX2_X1 port map( A => n9172, B => n2794, S => n1786, Z => n6363);
   U7403 : MUX2_X1 port map( A => n9173, B => n2783, S => n1786, Z => n6364);
   U7404 : MUX2_X1 port map( A => n9174, B => n2772, S => n1786, Z => n6365);
   U7405 : MUX2_X1 port map( A => n9175, B => n2761, S => n1786, Z => n6366);
   U7406 : MUX2_X1 port map( A => n9176, B => n2750, S => n1786, Z => n6367);
   U7407 : MUX2_X1 port map( A => n9177, B => n2739, S => n1786, Z => n6368);
   U7408 : MUX2_X1 port map( A => n9178, B => n2728, S => n1786, Z => n6369);
   U7409 : MUX2_X1 port map( A => n9179, B => n2717, S => n1786, Z => n6370);
   U7410 : MUX2_X1 port map( A => n9180, B => n2706, S => n1786, Z => n6371);
   U7411 : MUX2_X1 port map( A => n9181, B => n2599, S => n1786, Z => n6372);
   U7412 : MUX2_X1 port map( A => n9182, B => n2588, S => n1787, Z => n6373);
   U7413 : MUX2_X1 port map( A => n9183, B => n2577, S => n1787, Z => n6374);
   U7414 : MUX2_X1 port map( A => n9184, B => n2566, S => n1787, Z => n6375);
   U7415 : MUX2_X1 port map( A => n9185, B => n2555, S => n1787, Z => n6376);
   U7416 : MUX2_X1 port map( A => n9186, B => n2544, S => n1787, Z => n6377);
   U7417 : MUX2_X1 port map( A => n9187, B => n1829, S => n1787, Z => n6378);
   U7418 : MUX2_X1 port map( A => n9188, B => n1818, S => n1787, Z => n6379);
   U7419 : MUX2_X1 port map( A => n9189, B => n1807, S => n1787, Z => n6380);
   U7420 : MUX2_X1 port map( A => n3393, B => n2954, S => n1788, Z => n6317);
   U7421 : MUX2_X1 port map( A => n3395, B => n2943, S => n1788, Z => n6318);
   U7422 : MUX2_X1 port map( A => n3396, B => n2932, S => n1788, Z => n6319);
   U7423 : MUX2_X1 port map( A => n3397, B => n2917, S => n1788, Z => n6320);
   U7424 : MUX2_X1 port map( A => n3399, B => n2905, S => n1788, Z => n6321);
   U7425 : MUX2_X1 port map( A => n3401, B => n2893, S => n1788, Z => n6322);
   U7426 : MUX2_X1 port map( A => n3402, B => n2882, S => n1788, Z => n6323);
   U7427 : MUX2_X1 port map( A => n3404, B => n2871, S => n1788, Z => n6324);
   U7428 : MUX2_X1 port map( A => n3407, B => n2860, S => n1788, Z => n6325);
   U7429 : MUX2_X1 port map( A => n3408, B => n2849, S => n1788, Z => n6326);
   U7430 : MUX2_X1 port map( A => n3410, B => n2838, S => n1788, Z => n6327);
   U7431 : MUX2_X1 port map( A => n3411, B => n2827, S => n1788, Z => n6328);
   U7432 : MUX2_X1 port map( A => n3412, B => n2816, S => n1789, Z => n6329);
   U7433 : MUX2_X1 port map( A => n3414, B => n2805, S => n1789, Z => n6330);
   U7434 : MUX2_X1 port map( A => n9140, B => n2794, S => n1789, Z => n6331);
   U7435 : MUX2_X1 port map( A => n9141, B => n2783, S => n1789, Z => n6332);
   U7436 : MUX2_X1 port map( A => n9142, B => n2772, S => n1789, Z => n6333);
   U7437 : MUX2_X1 port map( A => n9143, B => n2761, S => n1789, Z => n6334);
   U7438 : MUX2_X1 port map( A => n9144, B => n2750, S => n1789, Z => n6335);
   U7439 : MUX2_X1 port map( A => n9145, B => n2739, S => n1789, Z => n6336);
   U7440 : MUX2_X1 port map( A => n9146, B => n2728, S => n1789, Z => n6337);
   U7441 : MUX2_X1 port map( A => n9147, B => n2717, S => n1789, Z => n6338);
   U7442 : MUX2_X1 port map( A => n9148, B => n2706, S => n1789, Z => n6339);
   U7443 : MUX2_X1 port map( A => n9149, B => n2599, S => n1789, Z => n6340);
   U7444 : MUX2_X1 port map( A => n9150, B => n2588, S => n1790, Z => n6341);
   U7445 : MUX2_X1 port map( A => n9151, B => n2577, S => n1790, Z => n6342);
   U7446 : MUX2_X1 port map( A => n9152, B => n2566, S => n1790, Z => n6343);
   U7447 : MUX2_X1 port map( A => n9153, B => n2555, S => n1790, Z => n6344);
   U7448 : MUX2_X1 port map( A => n9154, B => n2544, S => n1790, Z => n6345);
   U7449 : MUX2_X1 port map( A => n9155, B => n1829, S => n1790, Z => n6346);
   U7450 : MUX2_X1 port map( A => n9156, B => n1818, S => n1790, Z => n6347);
   U7451 : MUX2_X1 port map( A => n9157, B => n1807, S => n1790, Z => n6348);

end SYN_bhv;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity IR_DECODE_NBIT32_opBIT6_regBIT5 is

   port( CLK : in std_logic;  IR_26 : in std_logic_vector (25 downto 0);  
         OPCODE : in std_logic_vector (5 downto 0);  is_signed : in std_logic; 
         RS1, RS2, RD : out std_logic_vector (4 downto 0);  IMMEDIATE : out 
         std_logic_vector (31 downto 0));

end IR_DECODE_NBIT32_opBIT6_regBIT5;

architecture SYN_BEHAV of IR_DECODE_NBIT32_opBIT6_regBIT5 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X2
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component sign_eval_N_in26_N_out32
      port( IR_out : in std_logic_vector (25 downto 0);  signed_val : in 
            std_logic;  Immediate : out std_logic_vector (31 downto 0));
   end component;
   
   component sign_eval_N_in16_N_out32
      port( IR_out : in std_logic_vector (15 downto 0);  signed_val : in 
            std_logic;  Immediate : out std_logic_vector (31 downto 0));
   end component;
   
   component sign_eval_N_in5_N_out32
      port( IR_out : in std_logic_vector (4 downto 0);  signed_val : in 
            std_logic;  Immediate : out std_logic_vector (31 downto 0));
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal X_Logic0_port, IMMEDIATE_16_31_port, IMMEDIATE_16_15_port, 
      IMMEDIATE_16_14_port, IMMEDIATE_16_13_port, IMMEDIATE_16_12_port, 
      IMMEDIATE_16_11_port, IMMEDIATE_16_10_port, IMMEDIATE_16_9_port, 
      IMMEDIATE_16_8_port, IMMEDIATE_16_7_port, IMMEDIATE_16_6_port, 
      IMMEDIATE_16_5_port, IMMEDIATE_16_4_port, IMMEDIATE_16_3_port, 
      IMMEDIATE_16_2_port, IMMEDIATE_16_1_port, IMMEDIATE_16_0_port, N143, N144
      , N145, N146, N147, net105089, net137935, n1, n2, n3, n4, n5, n6, n7, n8,
      n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23,
      n_2212, n_2213, n_2214, n_2215, n_2216, n_2217, n_2218, n_2219, n_2220, 
      n_2221, n_2222, n_2223, n_2224, n_2225, n_2226, n_2227, n_2228, n_2229, 
      n_2230, n_2231, n_2232, n_2233, n_2234, n_2235, n_2236, n_2237, n_2238, 
      n_2239, n_2240, n_2241, n_2242, n_2243, n_2244, n_2245, n_2246, n_2247, 
      n_2248, n_2249, n_2250, n_2251, n_2252, n_2253, n_2254, n_2255, n_2256, 
      n_2257, n_2258, n_2259, n_2260, n_2261, n_2262, n_2263, n_2264, n_2265, 
      n_2266, n_2267, n_2268, n_2269, n_2270, n_2271, n_2272, n_2273, n_2274, 
      n_2275, n_2276, n_2277, n_2278, n_2279, n_2280, n_2281, n_2282, n_2283, 
      n_2284, n_2285, n_2286, n_2287, n_2288, n_2289, n_2290 : std_logic;

begin
   
   X_Logic0_port <= '0';
   RD_reg_4_inst : DLH_X1 port map( G => CLK, D => N147, Q => RD(4));
   RD_reg_3_inst : DLH_X1 port map( G => CLK, D => N146, Q => RD(3));
   RD_reg_2_inst : DLH_X1 port map( G => CLK, D => N145, Q => RD(2));
   RD_reg_1_inst : DLH_X1 port map( G => CLK, D => N144, Q => RD(1));
   RD_reg_0_inst : DLH_X1 port map( G => CLK, D => N143, Q => RD(0));
   IMMEDIATE_reg_31_inst : DLH_X1 port map( G => CLK, D => n7, Q => 
                           IMMEDIATE(31));
   IMMEDIATE_reg_30_inst : DLH_X1 port map( G => CLK, D => n23, Q => 
                           IMMEDIATE(30));
   IMMEDIATE_reg_29_inst : DLH_X1 port map( G => CLK, D => n23, Q => 
                           IMMEDIATE(29));
   IMMEDIATE_reg_28_inst : DLH_X1 port map( G => CLK, D => n7, Q => 
                           IMMEDIATE(28));
   IMMEDIATE_reg_27_inst : DLH_X1 port map( G => CLK, D => n7, Q => 
                           IMMEDIATE(27));
   IMMEDIATE_reg_26_inst : DLH_X1 port map( G => CLK, D => n23, Q => 
                           IMMEDIATE(26));
   IMMEDIATE_reg_25_inst : DLH_X1 port map( G => CLK, D => n23, Q => 
                           IMMEDIATE(25));
   IMMEDIATE_reg_24_inst : DLH_X1 port map( G => CLK, D => n7, Q => 
                           IMMEDIATE(24));
   IMMEDIATE_reg_23_inst : DLH_X1 port map( G => CLK, D => n7, Q => 
                           IMMEDIATE(23));
   IMMEDIATE_reg_22_inst : DLH_X1 port map( G => CLK, D => n23, Q => 
                           IMMEDIATE(22));
   IMMEDIATE_reg_21_inst : DLH_X1 port map( G => CLK, D => n23, Q => 
                           IMMEDIATE(21));
   IMMEDIATE_reg_20_inst : DLH_X1 port map( G => CLK, D => n7, Q => 
                           IMMEDIATE(20));
   IMMEDIATE_reg_19_inst : DLH_X1 port map( G => CLK, D => n7, Q => 
                           IMMEDIATE(19));
   IMMEDIATE_reg_18_inst : DLH_X1 port map( G => CLK, D => n23, Q => 
                           IMMEDIATE(18));
   IMMEDIATE_reg_17_inst : DLH_X1 port map( G => CLK, D => n23, Q => 
                           IMMEDIATE(17));
   IMMEDIATE_reg_16_inst : DLH_X1 port map( G => CLK, D => n7, Q => 
                           IMMEDIATE(16));
   IMMEDIATE_reg_15_inst : DLH_X1 port map( G => CLK, D => n22, Q => 
                           IMMEDIATE(15));
   IMMEDIATE_reg_14_inst : DLH_X1 port map( G => CLK, D => n21, Q => 
                           IMMEDIATE(14));
   IMMEDIATE_reg_13_inst : DLH_X1 port map( G => CLK, D => n20, Q => 
                           IMMEDIATE(13));
   IMMEDIATE_reg_12_inst : DLH_X1 port map( G => CLK, D => net105089, Q => 
                           IMMEDIATE(12));
   IMMEDIATE_reg_11_inst : DLH_X1 port map( G => CLK, D => n19, Q => 
                           IMMEDIATE(11));
   IMMEDIATE_reg_10_inst : DLH_X1 port map( G => CLK, D => n18, Q => 
                           IMMEDIATE(10));
   IMMEDIATE_reg_9_inst : DLH_X1 port map( G => CLK, D => n17, Q => 
                           IMMEDIATE(9));
   IMMEDIATE_reg_8_inst : DLH_X1 port map( G => CLK, D => n16, Q => 
                           IMMEDIATE(8));
   IMMEDIATE_reg_7_inst : DLH_X1 port map( G => CLK, D => n15, Q => 
                           IMMEDIATE(7));
   IMMEDIATE_reg_6_inst : DLH_X1 port map( G => CLK, D => n14, Q => 
                           IMMEDIATE(6));
   IMMEDIATE_reg_5_inst : DLH_X1 port map( G => CLK, D => n13, Q => 
                           IMMEDIATE(5));
   IMMEDIATE_reg_4_inst : DLH_X1 port map( G => CLK, D => n12, Q => 
                           IMMEDIATE(4));
   IMMEDIATE_reg_3_inst : DLH_X1 port map( G => CLK, D => n11, Q => 
                           IMMEDIATE(3));
   IMMEDIATE_reg_2_inst : DLH_X1 port map( G => CLK, D => n10, Q => 
                           IMMEDIATE(2));
   IMMEDIATE_reg_1_inst : DLH_X1 port map( G => CLK, D => n9, Q => IMMEDIATE(1)
                           );
   IMMEDIATE_reg_0_inst : DLH_X1 port map( G => CLK, D => n8, Q => IMMEDIATE(0)
                           );
   RS1_reg_4_inst : DLH_X1 port map( G => CLK, D => IR_26(25), Q => RS1(4));
   RS1_reg_3_inst : DLH_X1 port map( G => CLK, D => IR_26(24), Q => RS1(3));
   RS1_reg_2_inst : DLH_X1 port map( G => CLK, D => IR_26(23), Q => RS1(2));
   RS1_reg_1_inst : DLH_X1 port map( G => CLK, D => IR_26(22), Q => RS1(1));
   RS1_reg_0_inst : DLH_X1 port map( G => CLK, D => IR_26(21), Q => RS1(0));
   RS2_reg_4_inst : DLH_X1 port map( G => CLK, D => IR_26(20), Q => RS2(4));
   RS2_reg_3_inst : DLH_X1 port map( G => CLK, D => IR_26(19), Q => RS2(3));
   RS2_reg_2_inst : DLH_X1 port map( G => CLK, D => IR_26(18), Q => RS2(2));
   RS2_reg_1_inst : DLH_X1 port map( G => CLK, D => IR_26(17), Q => RS2(1));
   RS2_reg_0_inst : DLH_X1 port map( G => CLK, D => IR_26(16), Q => RS2(0));
   SIGN_EXTENSION_imm5 : sign_eval_N_in5_N_out32 port map( IR_out(4) => 
                           IR_26(15), IR_out(3) => IR_26(14), IR_out(2) => 
                           IR_26(13), IR_out(1) => IR_26(12), IR_out(0) => 
                           IR_26(11), signed_val => is_signed, Immediate(31) =>
                           n_2212, Immediate(30) => n_2213, Immediate(29) => 
                           n_2214, Immediate(28) => n_2215, Immediate(27) => 
                           n_2216, Immediate(26) => n_2217, Immediate(25) => 
                           n_2218, Immediate(24) => n_2219, Immediate(23) => 
                           n_2220, Immediate(22) => n_2221, Immediate(21) => 
                           n_2222, Immediate(20) => n_2223, Immediate(19) => 
                           n_2224, Immediate(18) => n_2225, Immediate(17) => 
                           n_2226, Immediate(16) => n_2227, Immediate(15) => 
                           n_2228, Immediate(14) => n_2229, Immediate(13) => 
                           n_2230, Immediate(12) => n_2231, Immediate(11) => 
                           n_2232, Immediate(10) => n_2233, Immediate(9) => 
                           n_2234, Immediate(8) => n_2235, Immediate(7) => 
                           n_2236, Immediate(6) => n_2237, Immediate(5) => 
                           n_2238, Immediate(4) => n_2239, Immediate(3) => 
                           n_2240, Immediate(2) => n_2241, Immediate(1) => 
                           n_2242, Immediate(0) => n_2243);
   SIGN_EXTENSION_imm16 : sign_eval_N_in16_N_out32 port map( IR_out(15) => 
                           IR_26(15), IR_out(14) => IR_26(14), IR_out(13) => 
                           IR_26(13), IR_out(12) => IR_26(12), IR_out(11) => 
                           IR_26(11), IR_out(10) => IR_26(10), IR_out(9) => 
                           IR_26(9), IR_out(8) => IR_26(8), IR_out(7) => 
                           IR_26(7), IR_out(6) => IR_26(6), IR_out(5) => 
                           IR_26(5), IR_out(4) => IR_26(4), IR_out(3) => 
                           IR_26(3), IR_out(2) => IR_26(2), IR_out(1) => 
                           IR_26(1), IR_out(0) => IR_26(0), signed_val => 
                           is_signed, Immediate(31) => IMMEDIATE_16_31_port, 
                           Immediate(30) => n_2244, Immediate(29) => n_2245, 
                           Immediate(28) => n_2246, Immediate(27) => n_2247, 
                           Immediate(26) => n_2248, Immediate(25) => n_2249, 
                           Immediate(24) => n_2250, Immediate(23) => n_2251, 
                           Immediate(22) => n_2252, Immediate(21) => n_2253, 
                           Immediate(20) => n_2254, Immediate(19) => n_2255, 
                           Immediate(18) => n_2256, Immediate(17) => n_2257, 
                           Immediate(16) => n_2258, Immediate(15) => 
                           IMMEDIATE_16_15_port, Immediate(14) => 
                           IMMEDIATE_16_14_port, Immediate(13) => 
                           IMMEDIATE_16_13_port, Immediate(12) => 
                           IMMEDIATE_16_12_port, Immediate(11) => 
                           IMMEDIATE_16_11_port, Immediate(10) => 
                           IMMEDIATE_16_10_port, Immediate(9) => 
                           IMMEDIATE_16_9_port, Immediate(8) => 
                           IMMEDIATE_16_8_port, Immediate(7) => 
                           IMMEDIATE_16_7_port, Immediate(6) => 
                           IMMEDIATE_16_6_port, Immediate(5) => 
                           IMMEDIATE_16_5_port, Immediate(4) => 
                           IMMEDIATE_16_4_port, Immediate(3) => 
                           IMMEDIATE_16_3_port, Immediate(2) => 
                           IMMEDIATE_16_2_port, Immediate(1) => 
                           IMMEDIATE_16_1_port, Immediate(0) => 
                           IMMEDIATE_16_0_port);
   SIGN_EXTENSION_imm26 : sign_eval_N_in26_N_out32 port map( IR_out(25) => 
                           IR_26(25), IR_out(24) => IR_26(24), IR_out(23) => 
                           IR_26(23), IR_out(22) => IR_26(22), IR_out(21) => 
                           IR_26(21), IR_out(20) => IR_26(20), IR_out(19) => 
                           IR_26(19), IR_out(18) => IR_26(18), IR_out(17) => 
                           IR_26(17), IR_out(16) => IR_26(16), IR_out(15) => 
                           IR_26(15), IR_out(14) => IR_26(14), IR_out(13) => 
                           IR_26(13), IR_out(12) => IR_26(12), IR_out(11) => 
                           IR_26(11), IR_out(10) => IR_26(10), IR_out(9) => 
                           IR_26(9), IR_out(8) => IR_26(8), IR_out(7) => 
                           IR_26(7), IR_out(6) => IR_26(6), IR_out(5) => 
                           IR_26(5), IR_out(4) => IR_26(4), IR_out(3) => 
                           IR_26(3), IR_out(2) => IR_26(2), IR_out(1) => 
                           IR_26(1), IR_out(0) => IR_26(0), signed_val => 
                           X_Logic0_port, Immediate(31) => n_2259, 
                           Immediate(30) => n_2260, Immediate(29) => n_2261, 
                           Immediate(28) => n_2262, Immediate(27) => n_2263, 
                           Immediate(26) => n_2264, Immediate(25) => n_2265, 
                           Immediate(24) => n_2266, Immediate(23) => n_2267, 
                           Immediate(22) => n_2268, Immediate(21) => n_2269, 
                           Immediate(20) => n_2270, Immediate(19) => n_2271, 
                           Immediate(18) => n_2272, Immediate(17) => n_2273, 
                           Immediate(16) => n_2274, Immediate(15) => n_2275, 
                           Immediate(14) => n_2276, Immediate(13) => n_2277, 
                           Immediate(12) => n_2278, Immediate(11) => n_2279, 
                           Immediate(10) => n_2280, Immediate(9) => n_2281, 
                           Immediate(8) => n_2282, Immediate(7) => n_2283, 
                           Immediate(6) => n_2284, Immediate(5) => n_2285, 
                           Immediate(4) => n_2286, Immediate(3) => n_2287, 
                           Immediate(2) => n_2288, Immediate(1) => n_2289, 
                           Immediate(0) => n_2290);
   U3 : NOR2_X1 port map( A1 => n1, A2 => n5, ZN => net105089);
   U4 : INV_X1 port map( A => IMMEDIATE_16_12_port, ZN => n5);
   U5 : AND2_X1 port map( A1 => n3, A2 => n2, ZN => n1);
   U6 : NOR3_X1 port map( A1 => OPCODE(2), A2 => OPCODE(1), A3 => OPCODE(0), ZN
                           => n2);
   U7 : NOR3_X1 port map( A1 => OPCODE(2), A2 => OPCODE(1), A3 => OPCODE(0), ZN
                           => n4);
   U8 : MUX2_X1 port map( A => IR_26(19), B => IR_26(14), S => n1, Z => N146);
   U9 : MUX2_X1 port map( A => IR_26(16), B => IR_26(11), S => n1, Z => N143);
   U10 : NOR3_X2 port map( A1 => OPCODE(5), A2 => OPCODE(4), A3 => OPCODE(3), 
                           ZN => n3);
   U11 : NAND2_X1 port map( A1 => n3, A2 => n4, ZN => net137935);
   U12 : NAND2_X1 port map( A1 => n3, A2 => n4, ZN => n6);
   U13 : AND2_X1 port map( A1 => IMMEDIATE_16_31_port, A2 => net137935, ZN => 
                           n7);
   U14 : AND2_X1 port map( A1 => IMMEDIATE_16_0_port, A2 => n6, ZN => n8);
   U15 : AND2_X1 port map( A1 => IMMEDIATE_16_1_port, A2 => n6, ZN => n9);
   U16 : AND2_X1 port map( A1 => IMMEDIATE_16_2_port, A2 => net137935, ZN => 
                           n10);
   U17 : AND2_X1 port map( A1 => IMMEDIATE_16_3_port, A2 => net137935, ZN => 
                           n11);
   U18 : AND2_X1 port map( A1 => IMMEDIATE_16_4_port, A2 => n6, ZN => n12);
   U19 : AND2_X1 port map( A1 => IMMEDIATE_16_5_port, A2 => n6, ZN => n13);
   U20 : AND2_X1 port map( A1 => IMMEDIATE_16_6_port, A2 => n6, ZN => n14);
   U21 : AND2_X1 port map( A1 => IMMEDIATE_16_7_port, A2 => n6, ZN => n15);
   U22 : AND2_X1 port map( A1 => IMMEDIATE_16_8_port, A2 => net137935, ZN => 
                           n16);
   U23 : AND2_X1 port map( A1 => IMMEDIATE_16_9_port, A2 => net137935, ZN => 
                           n17);
   U24 : AND2_X1 port map( A1 => IMMEDIATE_16_10_port, A2 => net137935, ZN => 
                           n18);
   U25 : AND2_X1 port map( A1 => IMMEDIATE_16_11_port, A2 => n6, ZN => n19);
   U26 : AND2_X1 port map( A1 => IMMEDIATE_16_13_port, A2 => net137935, ZN => 
                           n20);
   U27 : AND2_X1 port map( A1 => IMMEDIATE_16_14_port, A2 => n6, ZN => n21);
   U28 : AND2_X1 port map( A1 => IMMEDIATE_16_15_port, A2 => n6, ZN => n22);
   U29 : AND2_X1 port map( A1 => IMMEDIATE_16_31_port, A2 => net137935, ZN => 
                           n23);
   U30 : MUX2_X1 port map( A => IR_26(15), B => IR_26(20), S => n6, Z => N147);
   U31 : MUX2_X1 port map( A => IR_26(13), B => IR_26(18), S => net137935, Z =>
                           N145);
   U32 : MUX2_X1 port map( A => IR_26(12), B => IR_26(17), S => n6, Z => N144);

end SYN_BEHAV;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX21_GENERIC_NBIT32_0 is

   port( A, B : in std_logic_vector (31 downto 0);  SEL : in std_logic;  Y : 
         out std_logic_vector (31 downto 0));

end MUX21_GENERIC_NBIT32_0;

architecture SYN_struct of MUX21_GENERIC_NBIT32_0 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component MUX21_225
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_226
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_227
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_228
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_229
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_230
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_231
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_232
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_233
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_234
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_235
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_236
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_237
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_238
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_239
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_240
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_241
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_242
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_243
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_244
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_245
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_246
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_247
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_248
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_249
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_250
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_251
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_252
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_253
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_254
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_255
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_0
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   signal n1, n2, n3 : std_logic;

begin
   
   gen1_0 : MUX21_0 port map( A => A(0), B => B(0), S => n3, Y => Y(0));
   gen1_1 : MUX21_255 port map( A => A(1), B => B(1), S => n1, Y => Y(1));
   gen1_2 : MUX21_254 port map( A => A(2), B => B(2), S => n1, Y => Y(2));
   gen1_3 : MUX21_253 port map( A => A(3), B => B(3), S => n1, Y => Y(3));
   gen1_4 : MUX21_252 port map( A => A(4), B => B(4), S => n1, Y => Y(4));
   gen1_5 : MUX21_251 port map( A => A(5), B => B(5), S => n1, Y => Y(5));
   gen1_6 : MUX21_250 port map( A => A(6), B => B(6), S => n1, Y => Y(6));
   gen1_7 : MUX21_249 port map( A => A(7), B => B(7), S => n1, Y => Y(7));
   gen1_8 : MUX21_248 port map( A => A(8), B => B(8), S => n1, Y => Y(8));
   gen1_9 : MUX21_247 port map( A => A(9), B => B(9), S => n1, Y => Y(9));
   gen1_10 : MUX21_246 port map( A => A(10), B => B(10), S => n1, Y => Y(10));
   gen1_11 : MUX21_245 port map( A => A(11), B => B(11), S => n1, Y => Y(11));
   gen1_12 : MUX21_244 port map( A => A(12), B => B(12), S => n1, Y => Y(12));
   gen1_13 : MUX21_243 port map( A => A(13), B => B(13), S => n2, Y => Y(13));
   gen1_14 : MUX21_242 port map( A => A(14), B => B(14), S => n2, Y => Y(14));
   gen1_15 : MUX21_241 port map( A => A(15), B => B(15), S => n2, Y => Y(15));
   gen1_16 : MUX21_240 port map( A => A(16), B => B(16), S => n2, Y => Y(16));
   gen1_17 : MUX21_239 port map( A => A(17), B => B(17), S => n2, Y => Y(17));
   gen1_18 : MUX21_238 port map( A => A(18), B => B(18), S => n2, Y => Y(18));
   gen1_19 : MUX21_237 port map( A => A(19), B => B(19), S => n2, Y => Y(19));
   gen1_20 : MUX21_236 port map( A => A(20), B => B(20), S => n2, Y => Y(20));
   gen1_21 : MUX21_235 port map( A => A(21), B => B(21), S => n2, Y => Y(21));
   gen1_22 : MUX21_234 port map( A => A(22), B => B(22), S => n2, Y => Y(22));
   gen1_23 : MUX21_233 port map( A => A(23), B => B(23), S => n2, Y => Y(23));
   gen1_24 : MUX21_232 port map( A => A(24), B => B(24), S => n2, Y => Y(24));
   gen1_25 : MUX21_231 port map( A => A(25), B => B(25), S => n3, Y => Y(25));
   gen1_26 : MUX21_230 port map( A => A(26), B => B(26), S => n3, Y => Y(26));
   gen1_27 : MUX21_229 port map( A => A(27), B => B(27), S => n3, Y => Y(27));
   gen1_28 : MUX21_228 port map( A => A(28), B => B(28), S => n3, Y => Y(28));
   gen1_29 : MUX21_227 port map( A => A(29), B => B(29), S => n3, Y => Y(29));
   gen1_30 : MUX21_226 port map( A => A(30), B => B(30), S => n3, Y => Y(30));
   gen1_31 : MUX21_225 port map( A => A(31), B => B(31), S => n3, Y => Y(31));
   U1 : BUF_X1 port map( A => SEL, Z => n1);
   U2 : BUF_X1 port map( A => SEL, Z => n2);
   U3 : BUF_X1 port map( A => SEL, Z => n3);

end SYN_struct;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity regFFD_NBIT32_0 is

   port( CK, RESET, ENABLE : in std_logic;  D : in std_logic_vector (31 downto 
         0);  Q : out std_logic_vector (31 downto 0));

end regFFD_NBIT32_0;

architecture SYN_ASYNCHBEHAV of regFFD_NBIT32_0 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      , n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, 
      n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45
      , n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, 
      n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74
      , n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, 
      n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99 : std_logic;

begin
   
   Q_reg_31_inst : DFFR_X1 port map( D => n96, CK => CK, RN => n99, Q => Q(31),
                           QN => n64);
   Q_reg_30_inst : DFFR_X1 port map( D => n95, CK => CK, RN => n99, Q => Q(30),
                           QN => n63);
   Q_reg_29_inst : DFFR_X1 port map( D => n94, CK => CK, RN => n99, Q => Q(29),
                           QN => n62);
   Q_reg_28_inst : DFFR_X1 port map( D => n93, CK => CK, RN => n99, Q => Q(28),
                           QN => n61);
   Q_reg_27_inst : DFFR_X1 port map( D => n92, CK => CK, RN => n99, Q => Q(27),
                           QN => n60);
   Q_reg_26_inst : DFFR_X1 port map( D => n91, CK => CK, RN => n99, Q => Q(26),
                           QN => n59);
   Q_reg_25_inst : DFFR_X1 port map( D => n90, CK => CK, RN => n99, Q => Q(25),
                           QN => n58);
   Q_reg_24_inst : DFFR_X1 port map( D => n89, CK => CK, RN => n99, Q => Q(24),
                           QN => n57);
   Q_reg_23_inst : DFFR_X1 port map( D => n88, CK => CK, RN => n98, Q => Q(23),
                           QN => n56);
   Q_reg_22_inst : DFFR_X1 port map( D => n87, CK => CK, RN => n98, Q => Q(22),
                           QN => n55);
   Q_reg_21_inst : DFFR_X1 port map( D => n86, CK => CK, RN => n98, Q => Q(21),
                           QN => n54);
   Q_reg_20_inst : DFFR_X1 port map( D => n85, CK => CK, RN => n98, Q => Q(20),
                           QN => n53);
   Q_reg_19_inst : DFFR_X1 port map( D => n84, CK => CK, RN => n98, Q => Q(19),
                           QN => n52);
   Q_reg_18_inst : DFFR_X1 port map( D => n83, CK => CK, RN => n98, Q => Q(18),
                           QN => n51);
   Q_reg_17_inst : DFFR_X1 port map( D => n82, CK => CK, RN => n98, Q => Q(17),
                           QN => n50);
   Q_reg_16_inst : DFFR_X1 port map( D => n81, CK => CK, RN => n98, Q => Q(16),
                           QN => n49);
   Q_reg_15_inst : DFFR_X1 port map( D => n80, CK => CK, RN => n98, Q => Q(15),
                           QN => n48);
   Q_reg_14_inst : DFFR_X1 port map( D => n79, CK => CK, RN => n98, Q => Q(14),
                           QN => n47);
   Q_reg_13_inst : DFFR_X1 port map( D => n78, CK => CK, RN => n98, Q => Q(13),
                           QN => n46);
   Q_reg_12_inst : DFFR_X1 port map( D => n77, CK => CK, RN => n98, Q => Q(12),
                           QN => n45);
   Q_reg_11_inst : DFFR_X1 port map( D => n76, CK => CK, RN => n97, Q => Q(11),
                           QN => n44);
   Q_reg_10_inst : DFFR_X1 port map( D => n75, CK => CK, RN => n97, Q => Q(10),
                           QN => n43);
   Q_reg_9_inst : DFFR_X1 port map( D => n74, CK => CK, RN => n97, Q => Q(9), 
                           QN => n42);
   Q_reg_8_inst : DFFR_X1 port map( D => n73, CK => CK, RN => n97, Q => Q(8), 
                           QN => n41);
   Q_reg_7_inst : DFFR_X1 port map( D => n72, CK => CK, RN => n97, Q => Q(7), 
                           QN => n40);
   Q_reg_6_inst : DFFR_X1 port map( D => n71, CK => CK, RN => n97, Q => Q(6), 
                           QN => n39);
   Q_reg_5_inst : DFFR_X1 port map( D => n70, CK => CK, RN => n97, Q => Q(5), 
                           QN => n38);
   Q_reg_4_inst : DFFR_X1 port map( D => n69, CK => CK, RN => n97, Q => Q(4), 
                           QN => n37);
   Q_reg_3_inst : DFFR_X1 port map( D => n68, CK => CK, RN => n97, Q => Q(3), 
                           QN => n36);
   Q_reg_2_inst : DFFR_X1 port map( D => n67, CK => CK, RN => n97, Q => Q(2), 
                           QN => n35);
   Q_reg_1_inst : DFFR_X1 port map( D => n66, CK => CK, RN => n97, Q => Q(1), 
                           QN => n34);
   Q_reg_0_inst : DFFR_X1 port map( D => n65, CK => CK, RN => n97, Q => Q(0), 
                           QN => n33);
   U2 : BUF_X1 port map( A => RESET, Z => n97);
   U3 : BUF_X1 port map( A => RESET, Z => n98);
   U4 : BUF_X1 port map( A => RESET, Z => n99);
   U5 : OAI21_X1 port map( B1 => n33, B2 => ENABLE, A => n1, ZN => n65);
   U6 : NAND2_X1 port map( A1 => ENABLE, A2 => D(0), ZN => n1);
   U7 : OAI21_X1 port map( B1 => n34, B2 => ENABLE, A => n2, ZN => n66);
   U8 : NAND2_X1 port map( A1 => D(1), A2 => ENABLE, ZN => n2);
   U9 : OAI21_X1 port map( B1 => n35, B2 => ENABLE, A => n3, ZN => n67);
   U10 : NAND2_X1 port map( A1 => D(2), A2 => ENABLE, ZN => n3);
   U11 : OAI21_X1 port map( B1 => n36, B2 => ENABLE, A => n4, ZN => n68);
   U12 : NAND2_X1 port map( A1 => D(3), A2 => ENABLE, ZN => n4);
   U13 : OAI21_X1 port map( B1 => n37, B2 => ENABLE, A => n5, ZN => n69);
   U14 : NAND2_X1 port map( A1 => D(4), A2 => ENABLE, ZN => n5);
   U15 : OAI21_X1 port map( B1 => n38, B2 => ENABLE, A => n6, ZN => n70);
   U16 : NAND2_X1 port map( A1 => D(5), A2 => ENABLE, ZN => n6);
   U17 : OAI21_X1 port map( B1 => n39, B2 => ENABLE, A => n7, ZN => n71);
   U18 : NAND2_X1 port map( A1 => D(6), A2 => ENABLE, ZN => n7);
   U19 : OAI21_X1 port map( B1 => n40, B2 => ENABLE, A => n8, ZN => n72);
   U20 : NAND2_X1 port map( A1 => D(7), A2 => ENABLE, ZN => n8);
   U21 : OAI21_X1 port map( B1 => n41, B2 => ENABLE, A => n9, ZN => n73);
   U22 : NAND2_X1 port map( A1 => D(8), A2 => ENABLE, ZN => n9);
   U23 : OAI21_X1 port map( B1 => n42, B2 => ENABLE, A => n10, ZN => n74);
   U24 : NAND2_X1 port map( A1 => D(9), A2 => ENABLE, ZN => n10);
   U25 : OAI21_X1 port map( B1 => n43, B2 => ENABLE, A => n11, ZN => n75);
   U26 : NAND2_X1 port map( A1 => D(10), A2 => ENABLE, ZN => n11);
   U27 : OAI21_X1 port map( B1 => n44, B2 => ENABLE, A => n12, ZN => n76);
   U28 : NAND2_X1 port map( A1 => D(11), A2 => ENABLE, ZN => n12);
   U29 : OAI21_X1 port map( B1 => n45, B2 => ENABLE, A => n13, ZN => n77);
   U30 : NAND2_X1 port map( A1 => D(12), A2 => ENABLE, ZN => n13);
   U31 : OAI21_X1 port map( B1 => n46, B2 => ENABLE, A => n14, ZN => n78);
   U32 : NAND2_X1 port map( A1 => D(13), A2 => ENABLE, ZN => n14);
   U33 : OAI21_X1 port map( B1 => n47, B2 => ENABLE, A => n15, ZN => n79);
   U34 : NAND2_X1 port map( A1 => D(14), A2 => ENABLE, ZN => n15);
   U35 : OAI21_X1 port map( B1 => n48, B2 => ENABLE, A => n16, ZN => n80);
   U36 : NAND2_X1 port map( A1 => D(15), A2 => ENABLE, ZN => n16);
   U37 : OAI21_X1 port map( B1 => n49, B2 => ENABLE, A => n17, ZN => n81);
   U38 : NAND2_X1 port map( A1 => D(16), A2 => ENABLE, ZN => n17);
   U39 : OAI21_X1 port map( B1 => n50, B2 => ENABLE, A => n18, ZN => n82);
   U40 : NAND2_X1 port map( A1 => D(17), A2 => ENABLE, ZN => n18);
   U41 : OAI21_X1 port map( B1 => n51, B2 => ENABLE, A => n19, ZN => n83);
   U42 : NAND2_X1 port map( A1 => D(18), A2 => ENABLE, ZN => n19);
   U43 : OAI21_X1 port map( B1 => n52, B2 => ENABLE, A => n20, ZN => n84);
   U44 : NAND2_X1 port map( A1 => D(19), A2 => ENABLE, ZN => n20);
   U45 : OAI21_X1 port map( B1 => n53, B2 => ENABLE, A => n21, ZN => n85);
   U46 : NAND2_X1 port map( A1 => D(20), A2 => ENABLE, ZN => n21);
   U47 : OAI21_X1 port map( B1 => n54, B2 => ENABLE, A => n22, ZN => n86);
   U48 : NAND2_X1 port map( A1 => D(21), A2 => ENABLE, ZN => n22);
   U49 : OAI21_X1 port map( B1 => n55, B2 => ENABLE, A => n23, ZN => n87);
   U50 : NAND2_X1 port map( A1 => D(22), A2 => ENABLE, ZN => n23);
   U51 : OAI21_X1 port map( B1 => n56, B2 => ENABLE, A => n24, ZN => n88);
   U52 : NAND2_X1 port map( A1 => D(23), A2 => ENABLE, ZN => n24);
   U53 : OAI21_X1 port map( B1 => n57, B2 => ENABLE, A => n25, ZN => n89);
   U54 : NAND2_X1 port map( A1 => D(24), A2 => ENABLE, ZN => n25);
   U55 : OAI21_X1 port map( B1 => n58, B2 => ENABLE, A => n26, ZN => n90);
   U56 : NAND2_X1 port map( A1 => D(25), A2 => ENABLE, ZN => n26);
   U57 : OAI21_X1 port map( B1 => n59, B2 => ENABLE, A => n27, ZN => n91);
   U58 : NAND2_X1 port map( A1 => D(26), A2 => ENABLE, ZN => n27);
   U59 : OAI21_X1 port map( B1 => n60, B2 => ENABLE, A => n28, ZN => n92);
   U60 : NAND2_X1 port map( A1 => D(27), A2 => ENABLE, ZN => n28);
   U61 : OAI21_X1 port map( B1 => n61, B2 => ENABLE, A => n29, ZN => n93);
   U62 : NAND2_X1 port map( A1 => D(28), A2 => ENABLE, ZN => n29);
   U63 : OAI21_X1 port map( B1 => n62, B2 => ENABLE, A => n30, ZN => n94);
   U64 : NAND2_X1 port map( A1 => D(29), A2 => ENABLE, ZN => n30);
   U65 : OAI21_X1 port map( B1 => n63, B2 => ENABLE, A => n31, ZN => n95);
   U66 : NAND2_X1 port map( A1 => D(30), A2 => ENABLE, ZN => n31);
   U67 : OAI21_X1 port map( B1 => n64, B2 => ENABLE, A => n32, ZN => n96);
   U68 : NAND2_X1 port map( A1 => D(31), A2 => ENABLE, ZN => n32);

end SYN_ASYNCHBEHAV;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity DATAPTH_NBIT32_REG_BIT5 is

   port( CLK, RST : in std_logic;  PC, IR : in std_logic_vector (31 downto 0); 
         PC_OUT : out std_logic_vector (31 downto 0);  NPC_LATCH_EN, 
         ir_LATCH_EN, signed_op, trap_cs, ret_cs, RF1, RF2, WF1, 
         regImm_LATCH_EN, S1, S2, EN2, lhi_sel, jump_en, branch_cond, sb_op, RM
         , WM, EN3, S3 : in std_logic;  instruction_alu : in std_logic_vector 
         (0 to 5);  DATA_MEM_ADDR, DATA_MEM_IN : out std_logic_vector (31 
         downto 0);  DATA_MEM_OUT : in std_logic_vector (31 downto 0);  
         DATA_MEM_ENABLE, DATA_MEM_RM, DATA_MEM_WM : out std_logic);

end DATAPTH_NBIT32_REG_BIT5;

architecture SYN_STRUCTURAL of DATAPTH_NBIT32_REG_BIT5 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component BUF_X2
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component DATAPTH_NBIT32_REG_BIT5_DW01_inc_0
      port( A : in std_logic_vector (31 downto 0);  SUM : out std_logic_vector 
            (31 downto 0));
   end component;
   
   component MUX21_GENERIC_NBIT32_1
      port( A, B : in std_logic_vector (31 downto 0);  SEL : in std_logic;  Y :
            out std_logic_vector (31 downto 0));
   end component;
   
   component MUX21_GENERIC_NBIT32_2
      port( A, B : in std_logic_vector (31 downto 0);  SEL : in std_logic;  Y :
            out std_logic_vector (31 downto 0));
   end component;
   
   component regFFD_NBIT32_1
      port( CK, RESET, ENABLE : in std_logic;  D : in std_logic_vector (31 
            downto 0);  Q : out std_logic_vector (31 downto 0));
   end component;
   
   component FF_1
      port( CLK, RESET, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component FF_2
      port( CLK, RESET, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component FF_3
      port( CLK, RESET, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component regFFD_NBIT5_1
      port( CK, RESET, ENABLE : in std_logic;  D : in std_logic_vector (4 
            downto 0);  Q : out std_logic_vector (4 downto 0));
   end component;
   
   component regFFD_NBIT32_2
      port( CK, RESET, ENABLE : in std_logic;  D : in std_logic_vector (31 
            downto 0);  Q : out std_logic_vector (31 downto 0));
   end component;
   
   component regFFD_NBIT32_3
      port( CK, RESET, ENABLE : in std_logic;  D : in std_logic_vector (31 
            downto 0);  Q : out std_logic_vector (31 downto 0));
   end component;
   
   component load_data
      port( data_in : in std_logic_vector (31 downto 0);  signed_val, load_op :
            in std_logic;  load_type : in std_logic_vector (1 downto 0);  
            data_out : out std_logic_vector (31 downto 0));
   end component;
   
   component MUX21_GENERIC_NBIT32_3
      port( A, B : in std_logic_vector (31 downto 0);  SEL : in std_logic;  Y :
            out std_logic_vector (31 downto 0));
   end component;
   
   component regFFD_NBIT6_1
      port( CK, RESET, ENABLE : in std_logic;  D : in std_logic_vector (5 
            downto 0);  Q : out std_logic_vector (5 downto 0));
   end component;
   
   component FF_4
      port( CLK, RESET, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component regFFD_NBIT5_2
      port( CK, RESET, ENABLE : in std_logic;  D : in std_logic_vector (4 
            downto 0);  Q : out std_logic_vector (4 downto 0));
   end component;
   
   component regFFD_NBIT32_4
      port( CK, RESET, ENABLE : in std_logic;  D : in std_logic_vector (31 
            downto 0);  Q : out std_logic_vector (31 downto 0));
   end component;
   
   component FF_5
      port( CLK, RESET, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component regFFD_NBIT32_5
      port( CK, RESET, ENABLE : in std_logic;  D : in std_logic_vector (31 
            downto 0);  Q : out std_logic_vector (31 downto 0));
   end component;
   
   component FF_6
      port( CLK, RESET, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component MUX21_GENERIC_NBIT32_4
      port( A, B : in std_logic_vector (31 downto 0);  SEL : in std_logic;  Y :
            out std_logic_vector (31 downto 0));
   end component;
   
   component COND_BT_NBIT32
      port( ZERO_BIT, OPCODE_0, branch_op : in std_logic;  con_sign : out 
            std_logic);
   end component;
   
   component zero_eval_NBIT32
      port( input : in std_logic_vector (31 downto 0);  res : out std_logic);
   end component;
   
   component ALU_N32
      port( CLK : in std_logic;  FUNC : in std_logic_vector (0 to 5);  DATA1, 
            DATA2 : in std_logic_vector (31 downto 0);  OUT_ALU : out 
            std_logic_vector (31 downto 0));
   end component;
   
   component MUX21_GENERIC_NBIT32_5
      port( A, B : in std_logic_vector (31 downto 0);  SEL : in std_logic;  Y :
            out std_logic_vector (31 downto 0));
   end component;
   
   component MUX21_GENERIC_NBIT32_6
      port( A, B : in std_logic_vector (31 downto 0);  SEL : in std_logic;  Y :
            out std_logic_vector (31 downto 0));
   end component;
   
   component regFFD_NBIT32_6
      port( CK, RESET, ENABLE : in std_logic;  D : in std_logic_vector (31 
            downto 0);  Q : out std_logic_vector (31 downto 0));
   end component;
   
   component regFFD_NBIT6_0
      port( CK, RESET, ENABLE : in std_logic;  D : in std_logic_vector (5 
            downto 0);  Q : out std_logic_vector (5 downto 0));
   end component;
   
   component FF_7
      port( CLK, RESET, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component regFFD_NBIT5_0
      port( CK, RESET, ENABLE : in std_logic;  D : in std_logic_vector (4 
            downto 0);  Q : out std_logic_vector (4 downto 0));
   end component;
   
   component regFFD_NBIT32_7
      port( CK, RESET, ENABLE : in std_logic;  D : in std_logic_vector (31 
            downto 0);  Q : out std_logic_vector (31 downto 0));
   end component;
   
   component regFFD_NBIT32_8
      port( CK, RESET, ENABLE : in std_logic;  D : in std_logic_vector (31 
            downto 0);  Q : out std_logic_vector (31 downto 0));
   end component;
   
   component regFFD_NBIT32_9
      port( CK, RESET, ENABLE : in std_logic;  D : in std_logic_vector (31 
            downto 0);  Q : out std_logic_vector (31 downto 0));
   end component;
   
   component regFFD_NBIT32_10
      port( CK, RESET, ENABLE : in std_logic;  D : in std_logic_vector (31 
            downto 0);  Q : out std_logic_vector (31 downto 0));
   end component;
   
   component FF_0
      port( CLK, RESET, EN, D : in std_logic;  Q : out std_logic);
   end component;
   
   component windRF_M8_N8_F5_NBIT32
      port( CLK, RESET, ENABLE, CALL, RETRN : in std_logic;  FILL, SPILL : out 
            std_logic;  BUSin : in std_logic_vector (31 downto 0);  BUSout : 
            out std_logic_vector (31 downto 0);  RD1, RD2, WR : in std_logic;  
            ADD_WR, ADD_RD1, ADD_RD2 : in std_logic_vector (4 downto 0);  
            DATAIN : in std_logic_vector (31 downto 0);  OUT1, OUT2 : out 
            std_logic_vector (31 downto 0);  wr_signal : in std_logic);
   end component;
   
   component IR_DECODE_NBIT32_opBIT6_regBIT5
      port( CLK : in std_logic;  IR_26 : in std_logic_vector (25 downto 0);  
            OPCODE : in std_logic_vector (5 downto 0);  is_signed : in 
            std_logic;  RS1, RS2, RD : out std_logic_vector (4 downto 0);  
            IMMEDIATE : out std_logic_vector (31 downto 0));
   end component;
   
   component regFFD_NBIT32_11
      port( CK, RESET, ENABLE : in std_logic;  D : in std_logic_vector (31 
            downto 0);  Q : out std_logic_vector (31 downto 0));
   end component;
   
   component regFFD_NBIT32_12
      port( CK, RESET, ENABLE : in std_logic;  D : in std_logic_vector (31 
            downto 0);  Q : out std_logic_vector (31 downto 0));
   end component;
   
   component regFFD_NBIT32_13
      port( CK, RESET, ENABLE : in std_logic;  D : in std_logic_vector (31 
            downto 0);  Q : out std_logic_vector (31 downto 0));
   end component;
   
   component regFFD_NBIT32_14
      port( CK, RESET, ENABLE : in std_logic;  D : in std_logic_vector (31 
            downto 0);  Q : out std_logic_vector (31 downto 0));
   end component;
   
   component regFFD_NBIT32_15
      port( CK, RESET, ENABLE : in std_logic;  D : in std_logic_vector (31 
            downto 0);  Q : out std_logic_vector (31 downto 0));
   end component;
   
   component regFFD_NBIT32_16
      port( CK, RESET, ENABLE : in std_logic;  D : in std_logic_vector (31 
            downto 0);  Q : out std_logic_vector (31 downto 0));
   end component;
   
   component MUX21_GENERIC_NBIT32_0
      port( A, B : in std_logic_vector (31 downto 0);  SEL : in std_logic;  Y :
            out std_logic_vector (31 downto 0));
   end component;
   
   component regFFD_NBIT32_17
      port( CK, RESET, ENABLE : in std_logic;  D : in std_logic_vector (31 
            downto 0);  Q : out std_logic_vector (31 downto 0));
   end component;
   
   component regFFD_NBIT32_18
      port( CK, RESET, ENABLE : in std_logic;  D : in std_logic_vector (31 
            downto 0);  Q : out std_logic_vector (31 downto 0));
   end component;
   
   component regFFD_NBIT32_0
      port( CK, RESET, ENABLE : in std_logic;  D : in std_logic_vector (31 
            downto 0);  Q : out std_logic_vector (31 downto 0));
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component OAI33_X1
      port( A1, A2, A3, B1, B2, B3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, PC_fetch0_31_port, PC_fetch0_30_port, 
      PC_fetch0_29_port, PC_fetch0_28_port, PC_fetch0_27_port, 
      PC_fetch0_26_port, PC_fetch0_25_port, PC_fetch0_24_port, 
      PC_fetch0_23_port, PC_fetch0_22_port, PC_fetch0_21_port, 
      PC_fetch0_20_port, PC_fetch0_19_port, PC_fetch0_18_port, 
      PC_fetch0_17_port, PC_fetch0_16_port, PC_fetch0_15_port, 
      PC_fetch0_14_port, PC_fetch0_13_port, PC_fetch0_12_port, 
      PC_fetch0_11_port, PC_fetch0_10_port, PC_fetch0_9_port, PC_fetch0_8_port,
      PC_fetch0_7_port, PC_fetch0_6_port, PC_fetch0_5_port, PC_fetch0_4_port, 
      PC_fetch0_3_port, PC_fetch0_2_port, PC_fetch0_1_port, PC_fetch0_0_port, 
      NPC_31_port, NPC_30_port, NPC_29_port, NPC_28_port, NPC_27_port, 
      NPC_26_port, NPC_25_port, NPC_24_port, NPC_23_port, NPC_22_port, 
      NPC_21_port, NPC_20_port, NPC_19_port, NPC_18_port, NPC_17_port, 
      NPC_16_port, NPC_15_port, NPC_14_port, NPC_13_port, NPC_12_port, 
      NPC_11_port, NPC_10_port, NPC_9_port, NPC_8_port, NPC_7_port, NPC_6_port,
      NPC_5_port, NPC_4_port, NPC_3_port, NPC_2_port, NPC_1_port, NPC_0_port, 
      NPC_fetch1_31_port, NPC_fetch1_30_port, NPC_fetch1_29_port, 
      NPC_fetch1_28_port, NPC_fetch1_27_port, NPC_fetch1_26_port, 
      NPC_fetch1_25_port, NPC_fetch1_24_port, NPC_fetch1_23_port, 
      NPC_fetch1_22_port, NPC_fetch1_21_port, NPC_fetch1_20_port, 
      NPC_fetch1_19_port, NPC_fetch1_18_port, NPC_fetch1_17_port, 
      NPC_fetch1_16_port, NPC_fetch1_15_port, NPC_fetch1_14_port, 
      NPC_fetch1_13_port, NPC_fetch1_12_port, NPC_fetch1_11_port, 
      NPC_fetch1_10_port, NPC_fetch1_9_port, NPC_fetch1_8_port, 
      NPC_fetch1_7_port, NPC_fetch1_6_port, NPC_fetch1_5_port, 
      NPC_fetch1_4_port, NPC_fetch1_3_port, NPC_fetch1_2_port, 
      NPC_fetch1_1_port, NPC_fetch1_0_port, PC_fetch1_31_port, 
      PC_fetch1_30_port, PC_fetch1_29_port, PC_fetch1_28_port, 
      PC_fetch1_27_port, PC_fetch1_26_port, PC_fetch1_25_port, 
      PC_fetch1_24_port, PC_fetch1_23_port, PC_fetch1_22_port, 
      PC_fetch1_21_port, PC_fetch1_20_port, PC_fetch1_19_port, 
      PC_fetch1_18_port, PC_fetch1_17_port, PC_fetch1_16_port, 
      PC_fetch1_15_port, PC_fetch1_14_port, PC_fetch1_13_port, 
      PC_fetch1_12_port, PC_fetch1_11_port, PC_fetch1_10_port, PC_fetch1_9_port
      , PC_fetch1_8_port, PC_fetch1_7_port, PC_fetch1_6_port, PC_fetch1_5_port,
      PC_fetch1_4_port, PC_fetch1_3_port, PC_fetch1_2_port, PC_fetch1_1_port, 
      PC_fetch1_0_port, PC_OUT_i_31_port, PC_OUT_i_30_port, PC_OUT_i_29_port, 
      PC_OUT_i_28_port, PC_OUT_i_27_port, PC_OUT_i_26_port, PC_OUT_i_25_port, 
      PC_OUT_i_24_port, PC_OUT_i_23_port, PC_OUT_i_22_port, PC_OUT_i_21_port, 
      PC_OUT_i_20_port, PC_OUT_i_19_port, PC_OUT_i_18_port, PC_OUT_i_17_port, 
      PC_OUT_i_16_port, PC_OUT_i_15_port, PC_OUT_i_14_port, PC_OUT_i_13_port, 
      PC_OUT_i_12_port, PC_OUT_i_11_port, PC_OUT_i_10_port, PC_OUT_i_9_port, 
      PC_OUT_i_8_port, PC_OUT_i_7_port, PC_OUT_i_6_port, PC_OUT_i_5_port, 
      PC_OUT_i_4_port, PC_OUT_i_3_port, PC_OUT_i_2_port, PC_OUT_i_1_port, 
      PC_OUT_i_0_port, sel_npc, NPC_fetch_31_port, NPC_fetch_30_port, 
      NPC_fetch_29_port, NPC_fetch_28_port, NPC_fetch_27_port, 
      NPC_fetch_26_port, NPC_fetch_25_port, NPC_fetch_24_port, 
      NPC_fetch_23_port, NPC_fetch_22_port, NPC_fetch_21_port, 
      NPC_fetch_20_port, NPC_fetch_19_port, NPC_fetch_18_port, 
      NPC_fetch_17_port, NPC_fetch_16_port, NPC_fetch_15_port, 
      NPC_fetch_14_port, NPC_fetch_13_port, NPC_fetch_12_port, 
      NPC_fetch_11_port, NPC_fetch_10_port, NPC_fetch_9_port, NPC_fetch_8_port,
      NPC_fetch_7_port, NPC_fetch_6_port, NPC_fetch_5_port, NPC_fetch_4_port, 
      NPC_fetch_3_port, NPC_fetch_2_port, NPC_fetch_1_port, NPC_fetch_0_port, 
      PC_fetch_31_port, PC_fetch_30_port, PC_fetch_29_port, PC_fetch_28_port, 
      PC_fetch_27_port, PC_fetch_26_port, PC_fetch_25_port, PC_fetch_24_port, 
      PC_fetch_23_port, PC_fetch_22_port, PC_fetch_21_port, PC_fetch_20_port, 
      PC_fetch_19_port, PC_fetch_18_port, PC_fetch_17_port, PC_fetch_16_port, 
      PC_fetch_15_port, PC_fetch_14_port, PC_fetch_13_port, PC_fetch_12_port, 
      PC_fetch_11_port, PC_fetch_10_port, PC_fetch_9_port, PC_fetch_8_port, 
      PC_fetch_7_port, PC_fetch_6_port, PC_fetch_5_port, PC_fetch_4_port, 
      PC_fetch_3_port, PC_fetch_2_port, PC_fetch_1_port, PC_fetch_0_port, 
      ir_fetch_31_port, ir_fetch_30_port, ir_fetch_29_port, ir_fetch_28_port, 
      ir_fetch_27_port, ir_fetch_26_port, ir_fetch_25_port, ir_fetch_24_port, 
      ir_fetch_23_port, ir_fetch_22_port, ir_fetch_21_port, ir_fetch_20_port, 
      ir_fetch_19_port, ir_fetch_18_port, ir_fetch_17_port, ir_fetch_16_port, 
      ir_fetch_15_port, ir_fetch_14_port, ir_fetch_13_port, ir_fetch_12_port, 
      ir_fetch_11_port, ir_fetch_10_port, ir_fetch_9_port, ir_fetch_8_port, 
      ir_fetch_7_port, ir_fetch_6_port, ir_fetch_5_port, ir_fetch_4_port, 
      ir_fetch_3_port, ir_fetch_2_port, ir_fetch_1_port, ir_fetch_0_port, 
      NPC_Dec_31_port, NPC_Dec_30_port, NPC_Dec_29_port, NPC_Dec_28_port, 
      NPC_Dec_27_port, NPC_Dec_26_port, NPC_Dec_25_port, NPC_Dec_24_port, 
      NPC_Dec_23_port, NPC_Dec_22_port, NPC_Dec_21_port, NPC_Dec_20_port, 
      NPC_Dec_19_port, NPC_Dec_18_port, NPC_Dec_17_port, NPC_Dec_16_port, 
      NPC_Dec_15_port, NPC_Dec_14_port, NPC_Dec_13_port, NPC_Dec_12_port, 
      NPC_Dec_11_port, NPC_Dec_10_port, NPC_Dec_9_port, NPC_Dec_8_port, 
      NPC_Dec_7_port, NPC_Dec_6_port, NPC_Dec_5_port, NPC_Dec_4_port, 
      NPC_Dec_3_port, NPC_Dec_2_port, NPC_Dec_1_port, NPC_Dec_0_port, 
      IR_Dec_31_port, IR_Dec_30_port, IR_Dec_29_port, IR_Dec_28_port, 
      IR_Dec_27_port, IR_Dec_26_port, IR_Dec_25_port, IR_Dec_24_port, 
      IR_Dec_23_port, IR_Dec_22_port, IR_Dec_21_port, IR_Dec_20_port, 
      IR_Dec_19_port, IR_Dec_18_port, IR_Dec_17_port, IR_Dec_16_port, 
      IR_Dec_15_port, IR_Dec_14_port, IR_Dec_13_port, IR_Dec_12_port, 
      IR_Dec_11_port, IR_Dec_10_port, IR_Dec_9_port, IR_Dec_8_port, 
      IR_Dec_7_port, IR_Dec_6_port, IR_Dec_5_port, IR_Dec_4_port, IR_Dec_3_port
      , IR_Dec_2_port, IR_Dec_1_port, IR_Dec_0_port, RS1_4_port, RS1_3_port, 
      RS1_2_port, RS1_1_port, RS1_0_port, RS2_4_port, RS2_3_port, RS2_2_port, 
      RS2_1_port, RS2_0_port, RD_4_port, RD_3_port, RD_2_port, RD_1_port, 
      RD_0_port, Imm_31_port, Imm_30_port, Imm_29_port, Imm_28_port, 
      Imm_27_port, Imm_26_port, Imm_25_port, Imm_24_port, Imm_23_port, 
      Imm_22_port, Imm_21_port, Imm_20_port, Imm_19_port, Imm_18_port, 
      Imm_17_port, Imm_16_port, Imm_15_port, Imm_14_port, Imm_13_port, 
      Imm_12_port, Imm_11_port, Imm_10_port, Imm_9_port, Imm_8_port, Imm_7_port
      , Imm_6_port, Imm_5_port, Imm_4_port, Imm_3_port, Imm_2_port, Imm_1_port,
      Imm_0_port, RD_wb_4_port, RD_wb_3_port, RD_wb_2_port, RD_wb_1_port, 
      RD_wb_0_port, OUT_wb_31_port, OUT_wb_30_port, OUT_wb_29_port, 
      OUT_wb_28_port, OUT_wb_27_port, OUT_wb_26_port, OUT_wb_25_port, 
      OUT_wb_24_port, OUT_wb_23_port, OUT_wb_22_port, OUT_wb_21_port, 
      OUT_wb_20_port, OUT_wb_19_port, OUT_wb_18_port, OUT_wb_17_port, 
      OUT_wb_16_port, OUT_wb_15_port, OUT_wb_14_port, OUT_wb_13_port, 
      OUT_wb_12_port, OUT_wb_11_port, OUT_wb_10_port, OUT_wb_9_port, 
      OUT_wb_8_port, OUT_wb_7_port, OUT_wb_6_port, OUT_wb_5_port, OUT_wb_4_port
      , OUT_wb_3_port, OUT_wb_2_port, OUT_wb_1_port, OUT_wb_0_port, 
      regA_31_port, regA_30_port, regA_29_port, regA_28_port, regA_27_port, 
      regA_26_port, regA_25_port, regA_24_port, regA_23_port, regA_22_port, 
      regA_21_port, regA_20_port, regA_19_port, regA_18_port, regA_17_port, 
      regA_16_port, regA_15_port, regA_14_port, regA_13_port, regA_12_port, 
      regA_11_port, regA_10_port, regA_9_port, regA_8_port, regA_7_port, 
      regA_6_port, regA_5_port, regA_4_port, regA_3_port, regA_2_port, 
      regA_1_port, regA_0_port, regB_31_port, regB_30_port, regB_29_port, 
      regB_28_port, regB_27_port, regB_26_port, regB_25_port, regB_24_port, 
      regB_23_port, regB_22_port, regB_21_port, regB_20_port, regB_19_port, 
      regB_18_port, regB_17_port, regB_16_port, regB_15_port, regB_14_port, 
      regB_13_port, regB_12_port, regB_11_port, regB_10_port, regB_9_port, 
      regB_8_port, regB_7_port, regB_6_port, regB_5_port, regB_4_port, 
      regB_3_port, regB_2_port, regB_1_port, regB_0_port, wr_signal_wb, 
      signed_op_ex, NPC_ex_31_port, NPC_ex_30_port, NPC_ex_29_port, 
      NPC_ex_28_port, NPC_ex_27_port, NPC_ex_26_port, NPC_ex_25_port, 
      NPC_ex_24_port, NPC_ex_23_port, NPC_ex_22_port, NPC_ex_21_port, 
      NPC_ex_20_port, NPC_ex_19_port, NPC_ex_18_port, NPC_ex_17_port, 
      NPC_ex_16_port, NPC_ex_15_port, NPC_ex_14_port, NPC_ex_13_port, 
      NPC_ex_12_port, NPC_ex_11_port, NPC_ex_10_port, NPC_ex_9_port, 
      NPC_ex_8_port, NPC_ex_7_port, NPC_ex_6_port, NPC_ex_5_port, NPC_ex_4_port
      , NPC_ex_3_port, NPC_ex_2_port, NPC_ex_1_port, NPC_ex_0_port, 
      regA_ex_31_port, regA_ex_30_port, regA_ex_29_port, regA_ex_28_port, 
      regA_ex_27_port, regA_ex_26_port, regA_ex_25_port, regA_ex_24_port, 
      regA_ex_23_port, regA_ex_22_port, regA_ex_21_port, regA_ex_20_port, 
      regA_ex_19_port, regA_ex_18_port, regA_ex_17_port, regA_ex_16_port, 
      regA_ex_15_port, regA_ex_14_port, regA_ex_13_port, regA_ex_12_port, 
      regA_ex_11_port, regA_ex_10_port, regA_ex_9_port, regA_ex_8_port, 
      regA_ex_7_port, regA_ex_6_port, regA_ex_5_port, regA_ex_4_port, 
      regA_ex_3_port, regA_ex_2_port, regA_ex_1_port, regA_ex_0_port, 
      regB_ex_31_port, regB_ex_30_port, regB_ex_29_port, regB_ex_28_port, 
      regB_ex_27_port, regB_ex_26_port, regB_ex_25_port, regB_ex_24_port, 
      regB_ex_23_port, regB_ex_22_port, regB_ex_21_port, regB_ex_20_port, 
      regB_ex_19_port, regB_ex_18_port, regB_ex_17_port, regB_ex_16_port, 
      regB_ex_15_port, regB_ex_14_port, regB_ex_13_port, regB_ex_12_port, 
      regB_ex_11_port, regB_ex_10_port, regB_ex_9_port, regB_ex_8_port, 
      regB_ex_7_port, regB_ex_6_port, regB_ex_5_port, regB_ex_4_port, 
      regB_ex_3_port, regB_ex_2_port, regB_ex_1_port, regB_ex_0_port, 
      Imm_ex_31_port, Imm_ex_30_port, Imm_ex_29_port, Imm_ex_28_port, 
      Imm_ex_27_port, Imm_ex_26_port, Imm_ex_25_port, Imm_ex_24_port, 
      Imm_ex_23_port, Imm_ex_22_port, Imm_ex_21_port, Imm_ex_20_port, 
      Imm_ex_19_port, Imm_ex_18_port, Imm_ex_17_port, Imm_ex_16_port, 
      Imm_ex_15_port, Imm_ex_14_port, Imm_ex_13_port, Imm_ex_12_port, 
      Imm_ex_11_port, Imm_ex_10_port, Imm_ex_9_port, Imm_ex_8_port, 
      Imm_ex_7_port, Imm_ex_6_port, Imm_ex_5_port, Imm_ex_4_port, Imm_ex_3_port
      , Imm_ex_2_port, Imm_ex_1_port, Imm_ex_0_port, RD_ex_4_port, RD_ex_3_port
      , RD_ex_2_port, RD_ex_1_port, RD_ex_0_port, wr_signal_exe, 
      IR_26_ex_5_port, IR_26_ex_4_port, IR_26_ex_3_port, IR_26_ex_2_port, 
      IR_26_ex_1_port, IR_26_ex_0_port, LHI_ex_31_port, LHI_ex_30_port, 
      LHI_ex_29_port, LHI_ex_28_port, LHI_ex_27_port, LHI_ex_26_port, 
      LHI_ex_25_port, LHI_ex_24_port, LHI_ex_23_port, LHI_ex_22_port, 
      LHI_ex_21_port, LHI_ex_20_port, LHI_ex_19_port, LHI_ex_18_port, 
      LHI_ex_17_port, LHI_ex_16_port, LHI_ex_15_port, LHI_ex_14_port, 
      LHI_ex_13_port, LHI_ex_12_port, LHI_ex_11_port, LHI_ex_10_port, 
      LHI_ex_9_port, LHI_ex_8_port, LHI_ex_7_port, LHI_ex_6_port, LHI_ex_5_port
      , LHI_ex_4_port, LHI_ex_3_port, LHI_ex_2_port, LHI_ex_1_port, 
      LHI_ex_0_port, input1_ALU_31_port, input1_ALU_30_port, input1_ALU_29_port
      , input1_ALU_28_port, input1_ALU_27_port, input1_ALU_26_port, 
      input1_ALU_25_port, input1_ALU_24_port, input1_ALU_23_port, 
      input1_ALU_22_port, input1_ALU_21_port, input1_ALU_20_port, 
      input1_ALU_19_port, input1_ALU_18_port, input1_ALU_17_port, 
      input1_ALU_16_port, input1_ALU_15_port, input1_ALU_14_port, 
      input1_ALU_13_port, input1_ALU_12_port, input1_ALU_11_port, 
      input1_ALU_10_port, input1_ALU_9_port, input1_ALU_8_port, 
      input1_ALU_7_port, input1_ALU_6_port, input1_ALU_5_port, 
      input1_ALU_4_port, input1_ALU_3_port, input1_ALU_2_port, 
      input1_ALU_1_port, input1_ALU_0_port, input2_ALU_31_port, 
      input2_ALU_30_port, input2_ALU_29_port, input2_ALU_28_port, 
      input2_ALU_27_port, input2_ALU_26_port, input2_ALU_25_port, 
      input2_ALU_24_port, input2_ALU_23_port, input2_ALU_22_port, 
      input2_ALU_21_port, input2_ALU_20_port, input2_ALU_19_port, 
      input2_ALU_18_port, input2_ALU_17_port, input2_ALU_16_port, 
      input2_ALU_15_port, input2_ALU_14_port, input2_ALU_13_port, 
      input2_ALU_12_port, input2_ALU_11_port, input2_ALU_10_port, 
      input2_ALU_9_port, input2_ALU_8_port, input2_ALU_7_port, 
      input2_ALU_6_port, input2_ALU_5_port, input2_ALU_4_port, 
      input2_ALU_3_port, input2_ALU_2_port, input2_ALU_1_port, 
      input2_ALU_0_port, ALU_out_31_port, ALU_out_30_port, ALU_out_29_port, 
      ALU_out_28_port, ALU_out_27_port, ALU_out_26_port, ALU_out_25_port, 
      ALU_out_24_port, ALU_out_23_port, ALU_out_22_port, ALU_out_21_port, 
      ALU_out_20_port, ALU_out_19_port, ALU_out_18_port, ALU_out_17_port, 
      ALU_out_16_port, ALU_out_15_port, ALU_out_14_port, ALU_out_13_port, 
      ALU_out_12_port, ALU_out_11_port, ALU_out_10_port, ALU_out_9_port, 
      ALU_out_8_port, ALU_out_7_port, ALU_out_6_port, ALU_out_5_port, 
      ALU_out_4_port, ALU_out_3_port, ALU_out_2_port, ALU_out_1_port, 
      ALU_out_0_port, is_zero, cond, ALU_ex_31_port, ALU_ex_30_port, 
      ALU_ex_29_port, ALU_ex_28_port, ALU_ex_27_port, ALU_ex_26_port, 
      ALU_ex_25_port, ALU_ex_24_port, ALU_ex_23_port, ALU_ex_22_port, 
      ALU_ex_21_port, ALU_ex_20_port, ALU_ex_19_port, ALU_ex_18_port, 
      ALU_ex_17_port, ALU_ex_16_port, ALU_ex_15_port, ALU_ex_14_port, 
      ALU_ex_13_port, ALU_ex_12_port, ALU_ex_11_port, ALU_ex_10_port, 
      ALU_ex_9_port, ALU_ex_8_port, ALU_ex_7_port, ALU_ex_6_port, ALU_ex_5_port
      , ALU_ex_4_port, ALU_ex_3_port, ALU_ex_2_port, ALU_ex_1_port, 
      ALU_ex_0_port, signed_op_mem, NPC_mem_31_port, NPC_mem_30_port, 
      NPC_mem_29_port, NPC_mem_28_port, NPC_mem_27_port, NPC_mem_26_port, 
      NPC_mem_25_port, NPC_mem_24_port, NPC_mem_23_port, NPC_mem_22_port, 
      NPC_mem_21_port, NPC_mem_20_port, NPC_mem_19_port, NPC_mem_18_port, 
      NPC_mem_17_port, NPC_mem_16_port, NPC_mem_15_port, NPC_mem_14_port, 
      NPC_mem_13_port, NPC_mem_12_port, NPC_mem_11_port, NPC_mem_10_port, 
      NPC_mem_9_port, NPC_mem_8_port, NPC_mem_7_port, NPC_mem_6_port, 
      NPC_mem_5_port, NPC_mem_4_port, NPC_mem_3_port, NPC_mem_2_port, 
      NPC_mem_1_port, NPC_mem_0_port, cond_mem, regB_mem_31_port, 
      regB_mem_30_port, regB_mem_29_port, regB_mem_28_port, regB_mem_27_port, 
      regB_mem_26_port, regB_mem_25_port, regB_mem_24_port, regB_mem_23_port, 
      regB_mem_22_port, regB_mem_21_port, regB_mem_20_port, regB_mem_19_port, 
      regB_mem_18_port, regB_mem_17_port, regB_mem_16_port, regB_mem_15_port, 
      regB_mem_14_port, regB_mem_13_port, regB_mem_12_port, regB_mem_11_port, 
      regB_mem_10_port, regB_mem_9_port, regB_mem_8_port, regB_mem_7_port, 
      regB_mem_6_port, regB_mem_5_port, regB_mem_4_port, regB_mem_3_port, 
      regB_mem_2_port, regB_mem_1_port, regB_mem_0_port, RD_mem_4_port, 
      RD_mem_3_port, RD_mem_2_port, RD_mem_1_port, RD_mem_0_port, wr_signal_mem
      , IR_26_mem_5_port, IR_26_mem_4_port, IR_26_mem_3_port, IR_26_mem_2_port,
      IR_26_mem_1_port, IR_26_mem_0_port, sel_saved_reg, N13, wr_signal_mem1, 
      LMD_out_31_port, LMD_out_30_port, LMD_out_29_port, LMD_out_28_port, 
      LMD_out_27_port, LMD_out_26_port, LMD_out_25_port, LMD_out_24_port, 
      LMD_out_23_port, LMD_out_22_port, LMD_out_21_port, LMD_out_20_port, 
      LMD_out_19_port, LMD_out_18_port, LMD_out_17_port, LMD_out_16_port, 
      LMD_out_15_port, LMD_out_14_port, LMD_out_13_port, LMD_out_12_port, 
      LMD_out_11_port, LMD_out_10_port, LMD_out_9_port, LMD_out_8_port, 
      LMD_out_7_port, LMD_out_6_port, LMD_out_5_port, LMD_out_4_port, 
      LMD_out_3_port, LMD_out_2_port, LMD_out_1_port, LMD_out_0_port, 
      ALU_wb_31_port, ALU_wb_30_port, ALU_wb_29_port, ALU_wb_28_port, 
      ALU_wb_27_port, ALU_wb_26_port, ALU_wb_25_port, ALU_wb_24_port, 
      ALU_wb_23_port, ALU_wb_22_port, ALU_wb_21_port, ALU_wb_20_port, 
      ALU_wb_19_port, ALU_wb_18_port, ALU_wb_17_port, ALU_wb_16_port, 
      ALU_wb_15_port, ALU_wb_14_port, ALU_wb_13_port, ALU_wb_12_port, 
      ALU_wb_11_port, ALU_wb_10_port, ALU_wb_9_port, ALU_wb_8_port, 
      ALU_wb_7_port, ALU_wb_6_port, ALU_wb_5_port, ALU_wb_4_port, ALU_wb_3_port
      , ALU_wb_2_port, ALU_wb_1_port, ALU_wb_0_port, LMD_wb_31_port, 
      LMD_wb_30_port, LMD_wb_29_port, LMD_wb_28_port, LMD_wb_27_port, 
      LMD_wb_26_port, LMD_wb_25_port, LMD_wb_24_port, LMD_wb_23_port, 
      LMD_wb_22_port, LMD_wb_21_port, LMD_wb_20_port, LMD_wb_19_port, 
      LMD_wb_18_port, LMD_wb_17_port, LMD_wb_16_port, LMD_wb_15_port, 
      LMD_wb_14_port, LMD_wb_13_port, LMD_wb_12_port, LMD_wb_11_port, 
      LMD_wb_10_port, LMD_wb_9_port, LMD_wb_8_port, LMD_wb_7_port, 
      LMD_wb_6_port, LMD_wb_5_port, LMD_wb_4_port, LMD_wb_3_port, LMD_wb_2_port
      , LMD_wb_1_port, LMD_wb_0_port, sel_saved_reg_wb, NPC_wb_31_port, 
      NPC_wb_30_port, NPC_wb_29_port, NPC_wb_28_port, NPC_wb_27_port, 
      NPC_wb_26_port, NPC_wb_25_port, NPC_wb_24_port, NPC_wb_23_port, 
      NPC_wb_22_port, NPC_wb_21_port, NPC_wb_20_port, NPC_wb_19_port, 
      NPC_wb_18_port, NPC_wb_17_port, NPC_wb_16_port, NPC_wb_15_port, 
      NPC_wb_14_port, NPC_wb_13_port, NPC_wb_12_port, NPC_wb_11_port, 
      NPC_wb_10_port, NPC_wb_9_port, NPC_wb_8_port, NPC_wb_7_port, 
      NPC_wb_6_port, NPC_wb_5_port, NPC_wb_4_port, NPC_wb_3_port, NPC_wb_2_port
      , NPC_wb_1_port, NPC_wb_0_port, OUT_data_31_port, OUT_data_30_port, 
      OUT_data_29_port, OUT_data_28_port, OUT_data_27_port, OUT_data_26_port, 
      OUT_data_25_port, OUT_data_24_port, OUT_data_23_port, OUT_data_22_port, 
      OUT_data_21_port, OUT_data_20_port, OUT_data_19_port, OUT_data_18_port, 
      OUT_data_17_port, OUT_data_16_port, OUT_data_15_port, OUT_data_14_port, 
      OUT_data_13_port, OUT_data_12_port, OUT_data_11_port, OUT_data_10_port, 
      OUT_data_9_port, OUT_data_8_port, OUT_data_7_port, OUT_data_6_port, 
      OUT_data_5_port, OUT_data_4_port, OUT_data_3_port, OUT_data_2_port, 
      OUT_data_1_port, OUT_data_0_port, n21, n22, n23, n24, n25, n26, n27, n28,
      n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43
      , n44, n45, n46, n47, n48, n49, n50, n51, n52, n1, n2, n3, n4, n5, n6, n7
      , n8, n9, n10, n11, n12, n13_port, n14, n15, n16, n57, n58, n59, n60, n61
      , n_2291, n_2292, n_2293, n_2294, n_2295, n_2296, n_2297, n_2298, n_2299,
      n_2300, n_2301, n_2302, n_2303, n_2304, n_2305, n_2306, n_2307, n_2308, 
      n_2309, n_2310, n_2311, n_2312, n_2313, n_2314, n_2315, n_2316, n_2317, 
      n_2318, n_2319, n_2320, n_2321, n_2322, n_2323, n_2324, n_2325, n_2326, 
      n_2327, n_2328, n_2329, n_2330, n_2331, n_2332, n_2333, n_2334, n_2335, 
      n_2336, n_2337, n_2338, n_2339, n_2340, n_2341, n_2342, n_2343, n_2344, 
      n_2345, n_2346, n_2347, n_2348, n_2349, n_2350, n_2351, n_2352, n_2353, 
      n_2354, n_2355, n_2356, n_2357 : std_logic;

begin
   DATA_MEM_RM <= RM;
   DATA_MEM_WM <= WM;
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   DATA_MEM_ADDR_reg_31_inst : DLH_X1 port map( G => n5, D => ALU_ex_31_port, Q
                           => DATA_MEM_ADDR(31));
   DATA_MEM_ADDR_reg_30_inst : DLH_X1 port map( G => n5, D => ALU_ex_30_port, Q
                           => DATA_MEM_ADDR(30));
   DATA_MEM_ADDR_reg_29_inst : DLH_X1 port map( G => n5, D => ALU_ex_29_port, Q
                           => DATA_MEM_ADDR(29));
   DATA_MEM_ADDR_reg_28_inst : DLH_X1 port map( G => n5, D => ALU_ex_28_port, Q
                           => DATA_MEM_ADDR(28));
   DATA_MEM_ADDR_reg_27_inst : DLH_X1 port map( G => n5, D => ALU_ex_27_port, Q
                           => DATA_MEM_ADDR(27));
   DATA_MEM_ADDR_reg_26_inst : DLH_X1 port map( G => n5, D => ALU_ex_26_port, Q
                           => DATA_MEM_ADDR(26));
   DATA_MEM_ADDR_reg_25_inst : DLH_X1 port map( G => n5, D => ALU_ex_25_port, Q
                           => DATA_MEM_ADDR(25));
   DATA_MEM_ADDR_reg_24_inst : DLH_X1 port map( G => n5, D => ALU_ex_24_port, Q
                           => DATA_MEM_ADDR(24));
   DATA_MEM_ADDR_reg_23_inst : DLH_X1 port map( G => n5, D => ALU_ex_23_port, Q
                           => DATA_MEM_ADDR(23));
   DATA_MEM_ADDR_reg_22_inst : DLH_X1 port map( G => n5, D => ALU_ex_22_port, Q
                           => DATA_MEM_ADDR(22));
   DATA_MEM_ADDR_reg_21_inst : DLH_X1 port map( G => n5, D => ALU_ex_21_port, Q
                           => DATA_MEM_ADDR(21));
   DATA_MEM_ADDR_reg_20_inst : DLH_X1 port map( G => n6, D => ALU_ex_20_port, Q
                           => DATA_MEM_ADDR(20));
   DATA_MEM_ADDR_reg_19_inst : DLH_X1 port map( G => n6, D => ALU_ex_19_port, Q
                           => DATA_MEM_ADDR(19));
   DATA_MEM_ADDR_reg_18_inst : DLH_X1 port map( G => n6, D => ALU_ex_18_port, Q
                           => DATA_MEM_ADDR(18));
   DATA_MEM_ADDR_reg_17_inst : DLH_X1 port map( G => n6, D => ALU_ex_17_port, Q
                           => DATA_MEM_ADDR(17));
   DATA_MEM_ADDR_reg_16_inst : DLH_X1 port map( G => n6, D => ALU_ex_16_port, Q
                           => DATA_MEM_ADDR(16));
   DATA_MEM_ADDR_reg_15_inst : DLH_X1 port map( G => n6, D => ALU_ex_15_port, Q
                           => DATA_MEM_ADDR(15));
   DATA_MEM_ADDR_reg_14_inst : DLH_X1 port map( G => n6, D => ALU_ex_14_port, Q
                           => DATA_MEM_ADDR(14));
   DATA_MEM_ADDR_reg_13_inst : DLH_X1 port map( G => n6, D => ALU_ex_13_port, Q
                           => DATA_MEM_ADDR(13));
   DATA_MEM_ADDR_reg_12_inst : DLH_X1 port map( G => n6, D => ALU_ex_12_port, Q
                           => DATA_MEM_ADDR(12));
   DATA_MEM_ADDR_reg_11_inst : DLH_X1 port map( G => n6, D => ALU_ex_11_port, Q
                           => DATA_MEM_ADDR(11));
   DATA_MEM_ADDR_reg_10_inst : DLH_X1 port map( G => n6, D => ALU_ex_10_port, Q
                           => DATA_MEM_ADDR(10));
   DATA_MEM_ADDR_reg_9_inst : DLH_X1 port map( G => n7, D => ALU_ex_9_port, Q 
                           => DATA_MEM_ADDR(9));
   DATA_MEM_ADDR_reg_8_inst : DLH_X1 port map( G => n7, D => ALU_ex_8_port, Q 
                           => DATA_MEM_ADDR(8));
   DATA_MEM_ADDR_reg_7_inst : DLH_X1 port map( G => n7, D => ALU_ex_7_port, Q 
                           => DATA_MEM_ADDR(7));
   DATA_MEM_ADDR_reg_6_inst : DLH_X1 port map( G => n7, D => ALU_ex_6_port, Q 
                           => DATA_MEM_ADDR(6));
   DATA_MEM_ADDR_reg_5_inst : DLH_X1 port map( G => n7, D => ALU_ex_5_port, Q 
                           => DATA_MEM_ADDR(5));
   DATA_MEM_ADDR_reg_4_inst : DLH_X1 port map( G => n7, D => ALU_ex_4_port, Q 
                           => DATA_MEM_ADDR(4));
   DATA_MEM_ADDR_reg_3_inst : DLH_X1 port map( G => n7, D => ALU_ex_3_port, Q 
                           => DATA_MEM_ADDR(3));
   DATA_MEM_ADDR_reg_2_inst : DLH_X1 port map( G => n7, D => ALU_ex_2_port, Q 
                           => DATA_MEM_ADDR(2));
   DATA_MEM_ADDR_reg_1_inst : DLH_X1 port map( G => n7, D => ALU_ex_1_port, Q 
                           => DATA_MEM_ADDR(1));
   DATA_MEM_ADDR_reg_0_inst : DLH_X1 port map( G => n7, D => ALU_ex_0_port, Q 
                           => DATA_MEM_ADDR(0));
   U80 : OAI33_X1 port map( A1 => n15, A2 => IR_Dec_31_port, A3 => n2, B1 => 
                           n24, B2 => n13_port, B3 => n25, ZN => n23);
   U81 : XOR2_X1 port map( A => IR_Dec_27_port, B => IR_Dec_26_port, Z => n25);
   U82 : NAND3_X1 port map( A1 => n16, A2 => n14, A3 => n2, ZN => n24);
   U83 : NAND3_X1 port map( A1 => instruction_alu(3), A2 => instruction_alu(4),
                           A3 => instruction_alu(1), ZN => n52);
   pipeline_PCING : regFFD_NBIT32_0 port map( CK => CLK, RESET => n9, ENABLE =>
                           X_Logic1_port, D(31) => PC(31), D(30) => PC(30), 
                           D(29) => PC(29), D(28) => PC(28), D(27) => PC(27), 
                           D(26) => PC(26), D(25) => PC(25), D(24) => PC(24), 
                           D(23) => PC(23), D(22) => PC(22), D(21) => PC(21), 
                           D(20) => PC(20), D(19) => PC(19), D(18) => PC(18), 
                           D(17) => PC(17), D(16) => PC(16), D(15) => PC(15), 
                           D(14) => PC(14), D(13) => PC(13), D(12) => PC(12), 
                           D(11) => PC(11), D(10) => PC(10), D(9) => PC(9), 
                           D(8) => PC(8), D(7) => PC(7), D(6) => PC(6), D(5) =>
                           PC(5), D(4) => PC(4), D(3) => PC(3), D(2) => PC(2), 
                           D(1) => PC(1), D(0) => PC(0), Q(31) => 
                           PC_fetch0_31_port, Q(30) => PC_fetch0_30_port, Q(29)
                           => PC_fetch0_29_port, Q(28) => PC_fetch0_28_port, 
                           Q(27) => PC_fetch0_27_port, Q(26) => 
                           PC_fetch0_26_port, Q(25) => PC_fetch0_25_port, Q(24)
                           => PC_fetch0_24_port, Q(23) => PC_fetch0_23_port, 
                           Q(22) => PC_fetch0_22_port, Q(21) => 
                           PC_fetch0_21_port, Q(20) => PC_fetch0_20_port, Q(19)
                           => PC_fetch0_19_port, Q(18) => PC_fetch0_18_port, 
                           Q(17) => PC_fetch0_17_port, Q(16) => 
                           PC_fetch0_16_port, Q(15) => PC_fetch0_15_port, Q(14)
                           => PC_fetch0_14_port, Q(13) => PC_fetch0_13_port, 
                           Q(12) => PC_fetch0_12_port, Q(11) => 
                           PC_fetch0_11_port, Q(10) => PC_fetch0_10_port, Q(9) 
                           => PC_fetch0_9_port, Q(8) => PC_fetch0_8_port, Q(7) 
                           => PC_fetch0_7_port, Q(6) => PC_fetch0_6_port, Q(5) 
                           => PC_fetch0_5_port, Q(4) => PC_fetch0_4_port, Q(3) 
                           => PC_fetch0_3_port, Q(2) => PC_fetch0_2_port, Q(1) 
                           => PC_fetch0_1_port, Q(0) => PC_fetch0_0_port);
   pipeline_fetch1_NPC : regFFD_NBIT32_18 port map( CK => CLK, RESET => n9, 
                           ENABLE => NPC_LATCH_EN, D(31) => NPC_31_port, D(30) 
                           => NPC_30_port, D(29) => NPC_29_port, D(28) => 
                           NPC_28_port, D(27) => NPC_27_port, D(26) => 
                           NPC_26_port, D(25) => NPC_25_port, D(24) => 
                           NPC_24_port, D(23) => NPC_23_port, D(22) => 
                           NPC_22_port, D(21) => NPC_21_port, D(20) => 
                           NPC_20_port, D(19) => NPC_19_port, D(18) => 
                           NPC_18_port, D(17) => NPC_17_port, D(16) => 
                           NPC_16_port, D(15) => NPC_15_port, D(14) => 
                           NPC_14_port, D(13) => NPC_13_port, D(12) => 
                           NPC_12_port, D(11) => NPC_11_port, D(10) => 
                           NPC_10_port, D(9) => NPC_9_port, D(8) => NPC_8_port,
                           D(7) => NPC_7_port, D(6) => NPC_6_port, D(5) => 
                           NPC_5_port, D(4) => NPC_4_port, D(3) => NPC_3_port, 
                           D(2) => NPC_2_port, D(1) => NPC_1_port, D(0) => 
                           NPC_0_port, Q(31) => NPC_fetch1_31_port, Q(30) => 
                           NPC_fetch1_30_port, Q(29) => NPC_fetch1_29_port, 
                           Q(28) => NPC_fetch1_28_port, Q(27) => 
                           NPC_fetch1_27_port, Q(26) => NPC_fetch1_26_port, 
                           Q(25) => NPC_fetch1_25_port, Q(24) => 
                           NPC_fetch1_24_port, Q(23) => NPC_fetch1_23_port, 
                           Q(22) => NPC_fetch1_22_port, Q(21) => 
                           NPC_fetch1_21_port, Q(20) => NPC_fetch1_20_port, 
                           Q(19) => NPC_fetch1_19_port, Q(18) => 
                           NPC_fetch1_18_port, Q(17) => NPC_fetch1_17_port, 
                           Q(16) => NPC_fetch1_16_port, Q(15) => 
                           NPC_fetch1_15_port, Q(14) => NPC_fetch1_14_port, 
                           Q(13) => NPC_fetch1_13_port, Q(12) => 
                           NPC_fetch1_12_port, Q(11) => NPC_fetch1_11_port, 
                           Q(10) => NPC_fetch1_10_port, Q(9) => 
                           NPC_fetch1_9_port, Q(8) => NPC_fetch1_8_port, Q(7) 
                           => NPC_fetch1_7_port, Q(6) => NPC_fetch1_6_port, 
                           Q(5) => NPC_fetch1_5_port, Q(4) => NPC_fetch1_4_port
                           , Q(3) => NPC_fetch1_3_port, Q(2) => 
                           NPC_fetch1_2_port, Q(1) => NPC_fetch1_1_port, Q(0) 
                           => NPC_fetch1_0_port);
   pipeline_fetch1_PC : regFFD_NBIT32_17 port map( CK => CLK, RESET => n9, 
                           ENABLE => ir_LATCH_EN, D(31) => PC_fetch0_31_port, 
                           D(30) => PC_fetch0_30_port, D(29) => 
                           PC_fetch0_29_port, D(28) => PC_fetch0_28_port, D(27)
                           => PC_fetch0_27_port, D(26) => PC_fetch0_26_port, 
                           D(25) => PC_fetch0_25_port, D(24) => 
                           PC_fetch0_24_port, D(23) => PC_fetch0_23_port, D(22)
                           => PC_fetch0_22_port, D(21) => PC_fetch0_21_port, 
                           D(20) => PC_fetch0_20_port, D(19) => 
                           PC_fetch0_19_port, D(18) => PC_fetch0_18_port, D(17)
                           => PC_fetch0_17_port, D(16) => PC_fetch0_16_port, 
                           D(15) => PC_fetch0_15_port, D(14) => 
                           PC_fetch0_14_port, D(13) => PC_fetch0_13_port, D(12)
                           => PC_fetch0_12_port, D(11) => PC_fetch0_11_port, 
                           D(10) => PC_fetch0_10_port, D(9) => PC_fetch0_9_port
                           , D(8) => PC_fetch0_8_port, D(7) => PC_fetch0_7_port
                           , D(6) => PC_fetch0_6_port, D(5) => PC_fetch0_5_port
                           , D(4) => PC_fetch0_4_port, D(3) => PC_fetch0_3_port
                           , D(2) => PC_fetch0_2_port, D(1) => PC_fetch0_1_port
                           , D(0) => PC_fetch0_0_port, Q(31) => 
                           PC_fetch1_31_port, Q(30) => PC_fetch1_30_port, Q(29)
                           => PC_fetch1_29_port, Q(28) => PC_fetch1_28_port, 
                           Q(27) => PC_fetch1_27_port, Q(26) => 
                           PC_fetch1_26_port, Q(25) => PC_fetch1_25_port, Q(24)
                           => PC_fetch1_24_port, Q(23) => PC_fetch1_23_port, 
                           Q(22) => PC_fetch1_22_port, Q(21) => 
                           PC_fetch1_21_port, Q(20) => PC_fetch1_20_port, Q(19)
                           => PC_fetch1_19_port, Q(18) => PC_fetch1_18_port, 
                           Q(17) => PC_fetch1_17_port, Q(16) => 
                           PC_fetch1_16_port, Q(15) => PC_fetch1_15_port, Q(14)
                           => PC_fetch1_14_port, Q(13) => PC_fetch1_13_port, 
                           Q(12) => PC_fetch1_12_port, Q(11) => 
                           PC_fetch1_11_port, Q(10) => PC_fetch1_10_port, Q(9) 
                           => PC_fetch1_9_port, Q(8) => PC_fetch1_8_port, Q(7) 
                           => PC_fetch1_7_port, Q(6) => PC_fetch1_6_port, Q(5) 
                           => PC_fetch1_5_port, Q(4) => PC_fetch1_4_port, Q(3) 
                           => PC_fetch1_3_port, Q(2) => PC_fetch1_2_port, Q(1) 
                           => PC_fetch1_1_port, Q(0) => PC_fetch1_0_port);
   MUX_PC1 : MUX21_GENERIC_NBIT32_0 port map( A(31) => PC_OUT_i_31_port, A(30) 
                           => PC_OUT_i_30_port, A(29) => PC_OUT_i_29_port, 
                           A(28) => PC_OUT_i_28_port, A(27) => PC_OUT_i_27_port
                           , A(26) => PC_OUT_i_26_port, A(25) => 
                           PC_OUT_i_25_port, A(24) => PC_OUT_i_24_port, A(23) 
                           => PC_OUT_i_23_port, A(22) => PC_OUT_i_22_port, 
                           A(21) => PC_OUT_i_21_port, A(20) => PC_OUT_i_20_port
                           , A(19) => PC_OUT_i_19_port, A(18) => 
                           PC_OUT_i_18_port, A(17) => PC_OUT_i_17_port, A(16) 
                           => PC_OUT_i_16_port, A(15) => PC_OUT_i_15_port, 
                           A(14) => PC_OUT_i_14_port, A(13) => PC_OUT_i_13_port
                           , A(12) => PC_OUT_i_12_port, A(11) => 
                           PC_OUT_i_11_port, A(10) => PC_OUT_i_10_port, A(9) =>
                           PC_OUT_i_9_port, A(8) => PC_OUT_i_8_port, A(7) => 
                           PC_OUT_i_7_port, A(6) => PC_OUT_i_6_port, A(5) => 
                           PC_OUT_i_5_port, A(4) => PC_OUT_i_4_port, A(3) => 
                           PC_OUT_i_3_port, A(2) => PC_OUT_i_2_port, A(1) => 
                           PC_OUT_i_1_port, A(0) => PC_OUT_i_0_port, B(31) => 
                           NPC_fetch1_31_port, B(30) => NPC_fetch1_30_port, 
                           B(29) => NPC_fetch1_29_port, B(28) => 
                           NPC_fetch1_28_port, B(27) => NPC_fetch1_27_port, 
                           B(26) => NPC_fetch1_26_port, B(25) => 
                           NPC_fetch1_25_port, B(24) => NPC_fetch1_24_port, 
                           B(23) => NPC_fetch1_23_port, B(22) => 
                           NPC_fetch1_22_port, B(21) => NPC_fetch1_21_port, 
                           B(20) => NPC_fetch1_20_port, B(19) => 
                           NPC_fetch1_19_port, B(18) => NPC_fetch1_18_port, 
                           B(17) => NPC_fetch1_17_port, B(16) => 
                           NPC_fetch1_16_port, B(15) => NPC_fetch1_15_port, 
                           B(14) => NPC_fetch1_14_port, B(13) => 
                           NPC_fetch1_13_port, B(12) => NPC_fetch1_12_port, 
                           B(11) => NPC_fetch1_11_port, B(10) => 
                           NPC_fetch1_10_port, B(9) => NPC_fetch1_9_port, B(8) 
                           => NPC_fetch1_8_port, B(7) => NPC_fetch1_7_port, 
                           B(6) => NPC_fetch1_6_port, B(5) => NPC_fetch1_5_port
                           , B(4) => NPC_fetch1_4_port, B(3) => 
                           NPC_fetch1_3_port, B(2) => NPC_fetch1_2_port, B(1) 
                           => NPC_fetch1_1_port, B(0) => NPC_fetch1_0_port, SEL
                           => sel_npc, Y(31) => PC_OUT(31), Y(30) => PC_OUT(30)
                           , Y(29) => PC_OUT(29), Y(28) => PC_OUT(28), Y(27) =>
                           PC_OUT(27), Y(26) => PC_OUT(26), Y(25) => PC_OUT(25)
                           , Y(24) => PC_OUT(24), Y(23) => PC_OUT(23), Y(22) =>
                           PC_OUT(22), Y(21) => PC_OUT(21), Y(20) => PC_OUT(20)
                           , Y(19) => PC_OUT(19), Y(18) => PC_OUT(18), Y(17) =>
                           PC_OUT(17), Y(16) => PC_OUT(16), Y(15) => PC_OUT(15)
                           , Y(14) => PC_OUT(14), Y(13) => PC_OUT(13), Y(12) =>
                           PC_OUT(12), Y(11) => PC_OUT(11), Y(10) => PC_OUT(10)
                           , Y(9) => PC_OUT(9), Y(8) => PC_OUT(8), Y(7) => 
                           PC_OUT(7), Y(6) => PC_OUT(6), Y(5) => PC_OUT(5), 
                           Y(4) => PC_OUT(4), Y(3) => PC_OUT(3), Y(2) => 
                           PC_OUT(2), Y(1) => PC_OUT(1), Y(0) => PC_OUT(0));
   pipeline_fetch_NPC : regFFD_NBIT32_16 port map( CK => CLK, RESET => n9, 
                           ENABLE => NPC_LATCH_EN, D(31) => NPC_fetch1_31_port,
                           D(30) => NPC_fetch1_30_port, D(29) => 
                           NPC_fetch1_29_port, D(28) => NPC_fetch1_28_port, 
                           D(27) => NPC_fetch1_27_port, D(26) => 
                           NPC_fetch1_26_port, D(25) => NPC_fetch1_25_port, 
                           D(24) => NPC_fetch1_24_port, D(23) => 
                           NPC_fetch1_23_port, D(22) => NPC_fetch1_22_port, 
                           D(21) => NPC_fetch1_21_port, D(20) => 
                           NPC_fetch1_20_port, D(19) => NPC_fetch1_19_port, 
                           D(18) => NPC_fetch1_18_port, D(17) => 
                           NPC_fetch1_17_port, D(16) => NPC_fetch1_16_port, 
                           D(15) => NPC_fetch1_15_port, D(14) => 
                           NPC_fetch1_14_port, D(13) => NPC_fetch1_13_port, 
                           D(12) => NPC_fetch1_12_port, D(11) => 
                           NPC_fetch1_11_port, D(10) => NPC_fetch1_10_port, 
                           D(9) => NPC_fetch1_9_port, D(8) => NPC_fetch1_8_port
                           , D(7) => NPC_fetch1_7_port, D(6) => 
                           NPC_fetch1_6_port, D(5) => NPC_fetch1_5_port, D(4) 
                           => NPC_fetch1_4_port, D(3) => NPC_fetch1_3_port, 
                           D(2) => NPC_fetch1_2_port, D(1) => NPC_fetch1_1_port
                           , D(0) => NPC_fetch1_0_port, Q(31) => 
                           NPC_fetch_31_port, Q(30) => NPC_fetch_30_port, Q(29)
                           => NPC_fetch_29_port, Q(28) => NPC_fetch_28_port, 
                           Q(27) => NPC_fetch_27_port, Q(26) => 
                           NPC_fetch_26_port, Q(25) => NPC_fetch_25_port, Q(24)
                           => NPC_fetch_24_port, Q(23) => NPC_fetch_23_port, 
                           Q(22) => NPC_fetch_22_port, Q(21) => 
                           NPC_fetch_21_port, Q(20) => NPC_fetch_20_port, Q(19)
                           => NPC_fetch_19_port, Q(18) => NPC_fetch_18_port, 
                           Q(17) => NPC_fetch_17_port, Q(16) => 
                           NPC_fetch_16_port, Q(15) => NPC_fetch_15_port, Q(14)
                           => NPC_fetch_14_port, Q(13) => NPC_fetch_13_port, 
                           Q(12) => NPC_fetch_12_port, Q(11) => 
                           NPC_fetch_11_port, Q(10) => NPC_fetch_10_port, Q(9) 
                           => NPC_fetch_9_port, Q(8) => NPC_fetch_8_port, Q(7) 
                           => NPC_fetch_7_port, Q(6) => NPC_fetch_6_port, Q(5) 
                           => NPC_fetch_5_port, Q(4) => NPC_fetch_4_port, Q(3) 
                           => NPC_fetch_3_port, Q(2) => NPC_fetch_2_port, Q(1) 
                           => NPC_fetch_1_port, Q(0) => NPC_fetch_0_port);
   pipeline_fetch_PC : regFFD_NBIT32_15 port map( CK => CLK, RESET => n9, 
                           ENABLE => ir_LATCH_EN, D(31) => PC_fetch1_31_port, 
                           D(30) => PC_fetch1_30_port, D(29) => 
                           PC_fetch1_29_port, D(28) => PC_fetch1_28_port, D(27)
                           => PC_fetch1_27_port, D(26) => PC_fetch1_26_port, 
                           D(25) => PC_fetch1_25_port, D(24) => 
                           PC_fetch1_24_port, D(23) => PC_fetch1_23_port, D(22)
                           => PC_fetch1_22_port, D(21) => PC_fetch1_21_port, 
                           D(20) => PC_fetch1_20_port, D(19) => 
                           PC_fetch1_19_port, D(18) => PC_fetch1_18_port, D(17)
                           => PC_fetch1_17_port, D(16) => PC_fetch1_16_port, 
                           D(15) => PC_fetch1_15_port, D(14) => 
                           PC_fetch1_14_port, D(13) => PC_fetch1_13_port, D(12)
                           => PC_fetch1_12_port, D(11) => PC_fetch1_11_port, 
                           D(10) => PC_fetch1_10_port, D(9) => PC_fetch1_9_port
                           , D(8) => PC_fetch1_8_port, D(7) => PC_fetch1_7_port
                           , D(6) => PC_fetch1_6_port, D(5) => PC_fetch1_5_port
                           , D(4) => PC_fetch1_4_port, D(3) => PC_fetch1_3_port
                           , D(2) => PC_fetch1_2_port, D(1) => PC_fetch1_1_port
                           , D(0) => PC_fetch1_0_port, Q(31) => 
                           PC_fetch_31_port, Q(30) => PC_fetch_30_port, Q(29) 
                           => PC_fetch_29_port, Q(28) => PC_fetch_28_port, 
                           Q(27) => PC_fetch_27_port, Q(26) => PC_fetch_26_port
                           , Q(25) => PC_fetch_25_port, Q(24) => 
                           PC_fetch_24_port, Q(23) => PC_fetch_23_port, Q(22) 
                           => PC_fetch_22_port, Q(21) => PC_fetch_21_port, 
                           Q(20) => PC_fetch_20_port, Q(19) => PC_fetch_19_port
                           , Q(18) => PC_fetch_18_port, Q(17) => 
                           PC_fetch_17_port, Q(16) => PC_fetch_16_port, Q(15) 
                           => PC_fetch_15_port, Q(14) => PC_fetch_14_port, 
                           Q(13) => PC_fetch_13_port, Q(12) => PC_fetch_12_port
                           , Q(11) => PC_fetch_11_port, Q(10) => 
                           PC_fetch_10_port, Q(9) => PC_fetch_9_port, Q(8) => 
                           PC_fetch_8_port, Q(7) => PC_fetch_7_port, Q(6) => 
                           PC_fetch_6_port, Q(5) => PC_fetch_5_port, Q(4) => 
                           PC_fetch_4_port, Q(3) => PC_fetch_3_port, Q(2) => 
                           PC_fetch_2_port, Q(1) => PC_fetch_1_port, Q(0) => 
                           PC_fetch_0_port);
   pipeline_fetch_ir : regFFD_NBIT32_14 port map( CK => CLK, RESET => n9, 
                           ENABLE => ir_LATCH_EN, D(31) => IR(31), D(30) => 
                           IR(30), D(29) => IR(29), D(28) => IR(28), D(27) => 
                           IR(27), D(26) => IR(26), D(25) => IR(25), D(24) => 
                           IR(24), D(23) => IR(23), D(22) => IR(22), D(21) => 
                           IR(21), D(20) => IR(20), D(19) => IR(19), D(18) => 
                           IR(18), D(17) => IR(17), D(16) => IR(16), D(15) => 
                           IR(15), D(14) => IR(14), D(13) => IR(13), D(12) => 
                           IR(12), D(11) => IR(11), D(10) => IR(10), D(9) => 
                           IR(9), D(8) => IR(8), D(7) => IR(7), D(6) => IR(6), 
                           D(5) => IR(5), D(4) => IR(4), D(3) => IR(3), D(2) =>
                           IR(2), D(1) => IR(1), D(0) => IR(0), Q(31) => 
                           ir_fetch_31_port, Q(30) => ir_fetch_30_port, Q(29) 
                           => ir_fetch_29_port, Q(28) => ir_fetch_28_port, 
                           Q(27) => ir_fetch_27_port, Q(26) => ir_fetch_26_port
                           , Q(25) => ir_fetch_25_port, Q(24) => 
                           ir_fetch_24_port, Q(23) => ir_fetch_23_port, Q(22) 
                           => ir_fetch_22_port, Q(21) => ir_fetch_21_port, 
                           Q(20) => ir_fetch_20_port, Q(19) => ir_fetch_19_port
                           , Q(18) => ir_fetch_18_port, Q(17) => 
                           ir_fetch_17_port, Q(16) => ir_fetch_16_port, Q(15) 
                           => ir_fetch_15_port, Q(14) => ir_fetch_14_port, 
                           Q(13) => ir_fetch_13_port, Q(12) => ir_fetch_12_port
                           , Q(11) => ir_fetch_11_port, Q(10) => 
                           ir_fetch_10_port, Q(9) => ir_fetch_9_port, Q(8) => 
                           ir_fetch_8_port, Q(7) => ir_fetch_7_port, Q(6) => 
                           ir_fetch_6_port, Q(5) => ir_fetch_5_port, Q(4) => 
                           ir_fetch_4_port, Q(3) => ir_fetch_3_port, Q(2) => 
                           ir_fetch_2_port, Q(1) => ir_fetch_1_port, Q(0) => 
                           ir_fetch_0_port);
   pipeline_newpc1 : regFFD_NBIT32_13 port map( CK => CLK, RESET => n9, ENABLE 
                           => NPC_LATCH_EN, D(31) => NPC_fetch_31_port, D(30) 
                           => NPC_fetch_30_port, D(29) => NPC_fetch_29_port, 
                           D(28) => NPC_fetch_28_port, D(27) => 
                           NPC_fetch_27_port, D(26) => NPC_fetch_26_port, D(25)
                           => NPC_fetch_25_port, D(24) => NPC_fetch_24_port, 
                           D(23) => NPC_fetch_23_port, D(22) => 
                           NPC_fetch_22_port, D(21) => NPC_fetch_21_port, D(20)
                           => NPC_fetch_20_port, D(19) => NPC_fetch_19_port, 
                           D(18) => NPC_fetch_18_port, D(17) => 
                           NPC_fetch_17_port, D(16) => NPC_fetch_16_port, D(15)
                           => NPC_fetch_15_port, D(14) => NPC_fetch_14_port, 
                           D(13) => NPC_fetch_13_port, D(12) => 
                           NPC_fetch_12_port, D(11) => NPC_fetch_11_port, D(10)
                           => NPC_fetch_10_port, D(9) => NPC_fetch_9_port, D(8)
                           => NPC_fetch_8_port, D(7) => NPC_fetch_7_port, D(6) 
                           => NPC_fetch_6_port, D(5) => NPC_fetch_5_port, D(4) 
                           => NPC_fetch_4_port, D(3) => NPC_fetch_3_port, D(2) 
                           => NPC_fetch_2_port, D(1) => NPC_fetch_1_port, D(0) 
                           => NPC_fetch_0_port, Q(31) => NPC_Dec_31_port, Q(30)
                           => NPC_Dec_30_port, Q(29) => NPC_Dec_29_port, Q(28) 
                           => NPC_Dec_28_port, Q(27) => NPC_Dec_27_port, Q(26) 
                           => NPC_Dec_26_port, Q(25) => NPC_Dec_25_port, Q(24) 
                           => NPC_Dec_24_port, Q(23) => NPC_Dec_23_port, Q(22) 
                           => NPC_Dec_22_port, Q(21) => NPC_Dec_21_port, Q(20) 
                           => NPC_Dec_20_port, Q(19) => NPC_Dec_19_port, Q(18) 
                           => NPC_Dec_18_port, Q(17) => NPC_Dec_17_port, Q(16) 
                           => NPC_Dec_16_port, Q(15) => NPC_Dec_15_port, Q(14) 
                           => NPC_Dec_14_port, Q(13) => NPC_Dec_13_port, Q(12) 
                           => NPC_Dec_12_port, Q(11) => NPC_Dec_11_port, Q(10) 
                           => NPC_Dec_10_port, Q(9) => NPC_Dec_9_port, Q(8) => 
                           NPC_Dec_8_port, Q(7) => NPC_Dec_7_port, Q(6) => 
                           NPC_Dec_6_port, Q(5) => NPC_Dec_5_port, Q(4) => 
                           NPC_Dec_4_port, Q(3) => NPC_Dec_3_port, Q(2) => 
                           NPC_Dec_2_port, Q(1) => NPC_Dec_1_port, Q(0) => 
                           NPC_Dec_0_port);
   pipeline_pc1 : regFFD_NBIT32_12 port map( CK => CLK, RESET => n9, ENABLE => 
                           ir_LATCH_EN, D(31) => PC_fetch_31_port, D(30) => 
                           PC_fetch_30_port, D(29) => PC_fetch_29_port, D(28) 
                           => PC_fetch_28_port, D(27) => PC_fetch_27_port, 
                           D(26) => PC_fetch_26_port, D(25) => PC_fetch_25_port
                           , D(24) => PC_fetch_24_port, D(23) => 
                           PC_fetch_23_port, D(22) => PC_fetch_22_port, D(21) 
                           => PC_fetch_21_port, D(20) => PC_fetch_20_port, 
                           D(19) => PC_fetch_19_port, D(18) => PC_fetch_18_port
                           , D(17) => PC_fetch_17_port, D(16) => 
                           PC_fetch_16_port, D(15) => PC_fetch_15_port, D(14) 
                           => PC_fetch_14_port, D(13) => PC_fetch_13_port, 
                           D(12) => PC_fetch_12_port, D(11) => PC_fetch_11_port
                           , D(10) => PC_fetch_10_port, D(9) => PC_fetch_9_port
                           , D(8) => PC_fetch_8_port, D(7) => PC_fetch_7_port, 
                           D(6) => PC_fetch_6_port, D(5) => PC_fetch_5_port, 
                           D(4) => PC_fetch_4_port, D(3) => PC_fetch_3_port, 
                           D(2) => PC_fetch_2_port, D(1) => PC_fetch_1_port, 
                           D(0) => PC_fetch_0_port, Q(31) => n_2291, Q(30) => 
                           n_2292, Q(29) => n_2293, Q(28) => n_2294, Q(27) => 
                           n_2295, Q(26) => n_2296, Q(25) => n_2297, Q(24) => 
                           n_2298, Q(23) => n_2299, Q(22) => n_2300, Q(21) => 
                           n_2301, Q(20) => n_2302, Q(19) => n_2303, Q(18) => 
                           n_2304, Q(17) => n_2305, Q(16) => n_2306, Q(15) => 
                           n_2307, Q(14) => n_2308, Q(13) => n_2309, Q(12) => 
                           n_2310, Q(11) => n_2311, Q(10) => n_2312, Q(9) => 
                           n_2313, Q(8) => n_2314, Q(7) => n_2315, Q(6) => 
                           n_2316, Q(5) => n_2317, Q(4) => n_2318, Q(3) => 
                           n_2319, Q(2) => n_2320, Q(1) => n_2321, Q(0) => 
                           n_2322);
   pipeline_IR1 : regFFD_NBIT32_11 port map( CK => CLK, RESET => n9, ENABLE => 
                           ir_LATCH_EN, D(31) => ir_fetch_31_port, D(30) => 
                           ir_fetch_30_port, D(29) => ir_fetch_29_port, D(28) 
                           => ir_fetch_28_port, D(27) => ir_fetch_27_port, 
                           D(26) => ir_fetch_26_port, D(25) => ir_fetch_25_port
                           , D(24) => ir_fetch_24_port, D(23) => 
                           ir_fetch_23_port, D(22) => ir_fetch_22_port, D(21) 
                           => ir_fetch_21_port, D(20) => ir_fetch_20_port, 
                           D(19) => ir_fetch_19_port, D(18) => ir_fetch_18_port
                           , D(17) => ir_fetch_17_port, D(16) => 
                           ir_fetch_16_port, D(15) => ir_fetch_15_port, D(14) 
                           => ir_fetch_14_port, D(13) => ir_fetch_13_port, 
                           D(12) => ir_fetch_12_port, D(11) => ir_fetch_11_port
                           , D(10) => ir_fetch_10_port, D(9) => ir_fetch_9_port
                           , D(8) => ir_fetch_8_port, D(7) => ir_fetch_7_port, 
                           D(6) => ir_fetch_6_port, D(5) => ir_fetch_5_port, 
                           D(4) => ir_fetch_4_port, D(3) => ir_fetch_3_port, 
                           D(2) => ir_fetch_2_port, D(1) => ir_fetch_1_port, 
                           D(0) => ir_fetch_0_port, Q(31) => IR_Dec_31_port, 
                           Q(30) => IR_Dec_30_port, Q(29) => IR_Dec_29_port, 
                           Q(28) => IR_Dec_28_port, Q(27) => IR_Dec_27_port, 
                           Q(26) => IR_Dec_26_port, Q(25) => IR_Dec_25_port, 
                           Q(24) => IR_Dec_24_port, Q(23) => IR_Dec_23_port, 
                           Q(22) => IR_Dec_22_port, Q(21) => IR_Dec_21_port, 
                           Q(20) => IR_Dec_20_port, Q(19) => IR_Dec_19_port, 
                           Q(18) => IR_Dec_18_port, Q(17) => IR_Dec_17_port, 
                           Q(16) => IR_Dec_16_port, Q(15) => IR_Dec_15_port, 
                           Q(14) => IR_Dec_14_port, Q(13) => IR_Dec_13_port, 
                           Q(12) => IR_Dec_12_port, Q(11) => IR_Dec_11_port, 
                           Q(10) => IR_Dec_10_port, Q(9) => IR_Dec_9_port, Q(8)
                           => IR_Dec_8_port, Q(7) => IR_Dec_7_port, Q(6) => 
                           IR_Dec_6_port, Q(5) => IR_Dec_5_port, Q(4) => 
                           IR_Dec_4_port, Q(3) => IR_Dec_3_port, Q(2) => 
                           IR_Dec_2_port, Q(1) => IR_Dec_1_port, Q(0) => 
                           IR_Dec_0_port);
   IR_OP : IR_DECODE_NBIT32_opBIT6_regBIT5 port map( CLK => CLK, IR_26(25) => 
                           IR_Dec_25_port, IR_26(24) => IR_Dec_24_port, 
                           IR_26(23) => IR_Dec_23_port, IR_26(22) => 
                           IR_Dec_22_port, IR_26(21) => IR_Dec_21_port, 
                           IR_26(20) => IR_Dec_20_port, IR_26(19) => 
                           IR_Dec_19_port, IR_26(18) => IR_Dec_18_port, 
                           IR_26(17) => IR_Dec_17_port, IR_26(16) => 
                           IR_Dec_16_port, IR_26(15) => IR_Dec_15_port, 
                           IR_26(14) => IR_Dec_14_port, IR_26(13) => 
                           IR_Dec_13_port, IR_26(12) => IR_Dec_12_port, 
                           IR_26(11) => IR_Dec_11_port, IR_26(10) => 
                           IR_Dec_10_port, IR_26(9) => IR_Dec_9_port, IR_26(8) 
                           => IR_Dec_8_port, IR_26(7) => IR_Dec_7_port, 
                           IR_26(6) => IR_Dec_6_port, IR_26(5) => IR_Dec_5_port
                           , IR_26(4) => IR_Dec_4_port, IR_26(3) => 
                           IR_Dec_3_port, IR_26(2) => IR_Dec_2_port, IR_26(1) 
                           => IR_Dec_1_port, IR_26(0) => IR_Dec_0_port, 
                           OPCODE(5) => IR_Dec_31_port, OPCODE(4) => 
                           IR_Dec_30_port, OPCODE(3) => IR_Dec_29_port, 
                           OPCODE(2) => IR_Dec_28_port, OPCODE(1) => 
                           IR_Dec_27_port, OPCODE(0) => IR_Dec_26_port, 
                           is_signed => signed_op, RS1(4) => RS1_4_port, RS1(3)
                           => RS1_3_port, RS1(2) => RS1_2_port, RS1(1) => 
                           RS1_1_port, RS1(0) => RS1_0_port, RS2(4) => 
                           RS2_4_port, RS2(3) => RS2_3_port, RS2(2) => 
                           RS2_2_port, RS2(1) => RS2_1_port, RS2(0) => 
                           RS2_0_port, RD(4) => RD_4_port, RD(3) => RD_3_port, 
                           RD(2) => RD_2_port, RD(1) => RD_1_port, RD(0) => 
                           RD_0_port, IMMEDIATE(31) => Imm_31_port, 
                           IMMEDIATE(30) => Imm_30_port, IMMEDIATE(29) => 
                           Imm_29_port, IMMEDIATE(28) => Imm_28_port, 
                           IMMEDIATE(27) => Imm_27_port, IMMEDIATE(26) => 
                           Imm_26_port, IMMEDIATE(25) => Imm_25_port, 
                           IMMEDIATE(24) => Imm_24_port, IMMEDIATE(23) => 
                           Imm_23_port, IMMEDIATE(22) => Imm_22_port, 
                           IMMEDIATE(21) => Imm_21_port, IMMEDIATE(20) => 
                           Imm_20_port, IMMEDIATE(19) => Imm_19_port, 
                           IMMEDIATE(18) => Imm_18_port, IMMEDIATE(17) => 
                           Imm_17_port, IMMEDIATE(16) => Imm_16_port, 
                           IMMEDIATE(15) => Imm_15_port, IMMEDIATE(14) => 
                           Imm_14_port, IMMEDIATE(13) => Imm_13_port, 
                           IMMEDIATE(12) => Imm_12_port, IMMEDIATE(11) => 
                           Imm_11_port, IMMEDIATE(10) => Imm_10_port, 
                           IMMEDIATE(9) => Imm_9_port, IMMEDIATE(8) => 
                           Imm_8_port, IMMEDIATE(7) => Imm_7_port, IMMEDIATE(6)
                           => Imm_6_port, IMMEDIATE(5) => Imm_5_port, 
                           IMMEDIATE(4) => Imm_4_port, IMMEDIATE(3) => 
                           Imm_3_port, IMMEDIATE(2) => Imm_2_port, IMMEDIATE(1)
                           => Imm_1_port, IMMEDIATE(0) => Imm_0_port);
   RF : windRF_M8_N8_F5_NBIT32 port map( CLK => CLK, RESET => n8, ENABLE => 
                           X_Logic1_port, CALL => trap_cs, RETRN => ret_cs, 
                           FILL => n_2323, SPILL => n_2324, BUSin(31) => 
                           X_Logic0_port, BUSin(30) => X_Logic0_port, BUSin(29)
                           => X_Logic0_port, BUSin(28) => X_Logic0_port, 
                           BUSin(27) => X_Logic0_port, BUSin(26) => 
                           X_Logic0_port, BUSin(25) => X_Logic0_port, BUSin(24)
                           => X_Logic0_port, BUSin(23) => X_Logic0_port, 
                           BUSin(22) => X_Logic0_port, BUSin(21) => 
                           X_Logic0_port, BUSin(20) => X_Logic0_port, BUSin(19)
                           => X_Logic0_port, BUSin(18) => X_Logic0_port, 
                           BUSin(17) => X_Logic0_port, BUSin(16) => 
                           X_Logic0_port, BUSin(15) => X_Logic0_port, BUSin(14)
                           => X_Logic0_port, BUSin(13) => X_Logic0_port, 
                           BUSin(12) => X_Logic0_port, BUSin(11) => 
                           X_Logic0_port, BUSin(10) => X_Logic0_port, BUSin(9) 
                           => X_Logic0_port, BUSin(8) => X_Logic0_port, 
                           BUSin(7) => X_Logic0_port, BUSin(6) => X_Logic0_port
                           , BUSin(5) => X_Logic0_port, BUSin(4) => 
                           X_Logic0_port, BUSin(3) => X_Logic0_port, BUSin(2) 
                           => X_Logic0_port, BUSin(1) => X_Logic0_port, 
                           BUSin(0) => X_Logic0_port, BUSout(31) => n_2325, 
                           BUSout(30) => n_2326, BUSout(29) => n_2327, 
                           BUSout(28) => n_2328, BUSout(27) => n_2329, 
                           BUSout(26) => n_2330, BUSout(25) => n_2331, 
                           BUSout(24) => n_2332, BUSout(23) => n_2333, 
                           BUSout(22) => n_2334, BUSout(21) => n_2335, 
                           BUSout(20) => n_2336, BUSout(19) => n_2337, 
                           BUSout(18) => n_2338, BUSout(17) => n_2339, 
                           BUSout(16) => n_2340, BUSout(15) => n_2341, 
                           BUSout(14) => n_2342, BUSout(13) => n_2343, 
                           BUSout(12) => n_2344, BUSout(11) => n_2345, 
                           BUSout(10) => n_2346, BUSout(9) => n_2347, BUSout(8)
                           => n_2348, BUSout(7) => n_2349, BUSout(6) => n_2350,
                           BUSout(5) => n_2351, BUSout(4) => n_2352, BUSout(3) 
                           => n_2353, BUSout(2) => n_2354, BUSout(1) => n_2355,
                           BUSout(0) => n_2356, RD1 => RF1, RD2 => RF2, WR => 
                           WF1, ADD_WR(4) => RD_wb_4_port, ADD_WR(3) => 
                           RD_wb_3_port, ADD_WR(2) => RD_wb_2_port, ADD_WR(1) 
                           => RD_wb_1_port, ADD_WR(0) => RD_wb_0_port, 
                           ADD_RD1(4) => RS1_4_port, ADD_RD1(3) => RS1_3_port, 
                           ADD_RD1(2) => RS1_2_port, ADD_RD1(1) => RS1_1_port, 
                           ADD_RD1(0) => RS1_0_port, ADD_RD2(4) => RS2_4_port, 
                           ADD_RD2(3) => RS2_3_port, ADD_RD2(2) => RS2_2_port, 
                           ADD_RD2(1) => RS2_1_port, ADD_RD2(0) => RS2_0_port, 
                           DATAIN(31) => OUT_wb_31_port, DATAIN(30) => 
                           OUT_wb_30_port, DATAIN(29) => OUT_wb_29_port, 
                           DATAIN(28) => OUT_wb_28_port, DATAIN(27) => 
                           OUT_wb_27_port, DATAIN(26) => OUT_wb_26_port, 
                           DATAIN(25) => OUT_wb_25_port, DATAIN(24) => 
                           OUT_wb_24_port, DATAIN(23) => OUT_wb_23_port, 
                           DATAIN(22) => OUT_wb_22_port, DATAIN(21) => 
                           OUT_wb_21_port, DATAIN(20) => OUT_wb_20_port, 
                           DATAIN(19) => OUT_wb_19_port, DATAIN(18) => 
                           OUT_wb_18_port, DATAIN(17) => OUT_wb_17_port, 
                           DATAIN(16) => OUT_wb_16_port, DATAIN(15) => 
                           OUT_wb_15_port, DATAIN(14) => OUT_wb_14_port, 
                           DATAIN(13) => OUT_wb_13_port, DATAIN(12) => 
                           OUT_wb_12_port, DATAIN(11) => OUT_wb_11_port, 
                           DATAIN(10) => OUT_wb_10_port, DATAIN(9) => 
                           OUT_wb_9_port, DATAIN(8) => OUT_wb_8_port, DATAIN(7)
                           => OUT_wb_7_port, DATAIN(6) => OUT_wb_6_port, 
                           DATAIN(5) => OUT_wb_5_port, DATAIN(4) => 
                           OUT_wb_4_port, DATAIN(3) => OUT_wb_3_port, DATAIN(2)
                           => OUT_wb_2_port, DATAIN(1) => OUT_wb_1_port, 
                           DATAIN(0) => OUT_wb_0_port, OUT1(31) => regA_31_port
                           , OUT1(30) => regA_30_port, OUT1(29) => regA_29_port
                           , OUT1(28) => regA_28_port, OUT1(27) => regA_27_port
                           , OUT1(26) => regA_26_port, OUT1(25) => regA_25_port
                           , OUT1(24) => regA_24_port, OUT1(23) => regA_23_port
                           , OUT1(22) => regA_22_port, OUT1(21) => regA_21_port
                           , OUT1(20) => regA_20_port, OUT1(19) => regA_19_port
                           , OUT1(18) => regA_18_port, OUT1(17) => regA_17_port
                           , OUT1(16) => regA_16_port, OUT1(15) => regA_15_port
                           , OUT1(14) => regA_14_port, OUT1(13) => regA_13_port
                           , OUT1(12) => regA_12_port, OUT1(11) => regA_11_port
                           , OUT1(10) => regA_10_port, OUT1(9) => regA_9_port, 
                           OUT1(8) => regA_8_port, OUT1(7) => regA_7_port, 
                           OUT1(6) => regA_6_port, OUT1(5) => regA_5_port, 
                           OUT1(4) => regA_4_port, OUT1(3) => regA_3_port, 
                           OUT1(2) => regA_2_port, OUT1(1) => regA_1_port, 
                           OUT1(0) => regA_0_port, OUT2(31) => regB_31_port, 
                           OUT2(30) => regB_30_port, OUT2(29) => regB_29_port, 
                           OUT2(28) => regB_28_port, OUT2(27) => regB_27_port, 
                           OUT2(26) => regB_26_port, OUT2(25) => regB_25_port, 
                           OUT2(24) => regB_24_port, OUT2(23) => regB_23_port, 
                           OUT2(22) => regB_22_port, OUT2(21) => regB_21_port, 
                           OUT2(20) => regB_20_port, OUT2(19) => regB_19_port, 
                           OUT2(18) => regB_18_port, OUT2(17) => regB_17_port, 
                           OUT2(16) => regB_16_port, OUT2(15) => regB_15_port, 
                           OUT2(14) => regB_14_port, OUT2(13) => regB_13_port, 
                           OUT2(12) => regB_12_port, OUT2(11) => regB_11_port, 
                           OUT2(10) => regB_10_port, OUT2(9) => regB_9_port, 
                           OUT2(8) => regB_8_port, OUT2(7) => regB_7_port, 
                           OUT2(6) => regB_6_port, OUT2(5) => regB_5_port, 
                           OUT2(4) => regB_4_port, OUT2(3) => regB_3_port, 
                           OUT2(2) => regB_2_port, OUT2(1) => regB_1_port, 
                           OUT2(0) => regB_0_port, wr_signal => wr_signal_wb);
   pipeline_sign2 : FF_0 port map( CLK => CLK, RESET => n9, EN => X_Logic1_port
                           , D => signed_op, Q => signed_op_ex);
   pipeline_newpc2 : regFFD_NBIT32_10 port map( CK => CLK, RESET => n9, ENABLE 
                           => X_Logic1_port, D(31) => NPC_Dec_31_port, D(30) =>
                           NPC_Dec_30_port, D(29) => NPC_Dec_29_port, D(28) => 
                           NPC_Dec_28_port, D(27) => NPC_Dec_27_port, D(26) => 
                           NPC_Dec_26_port, D(25) => NPC_Dec_25_port, D(24) => 
                           NPC_Dec_24_port, D(23) => NPC_Dec_23_port, D(22) => 
                           NPC_Dec_22_port, D(21) => NPC_Dec_21_port, D(20) => 
                           NPC_Dec_20_port, D(19) => NPC_Dec_19_port, D(18) => 
                           NPC_Dec_18_port, D(17) => NPC_Dec_17_port, D(16) => 
                           NPC_Dec_16_port, D(15) => NPC_Dec_15_port, D(14) => 
                           NPC_Dec_14_port, D(13) => NPC_Dec_13_port, D(12) => 
                           NPC_Dec_12_port, D(11) => NPC_Dec_11_port, D(10) => 
                           NPC_Dec_10_port, D(9) => NPC_Dec_9_port, D(8) => 
                           NPC_Dec_8_port, D(7) => NPC_Dec_7_port, D(6) => 
                           NPC_Dec_6_port, D(5) => NPC_Dec_5_port, D(4) => 
                           NPC_Dec_4_port, D(3) => NPC_Dec_3_port, D(2) => 
                           NPC_Dec_2_port, D(1) => NPC_Dec_1_port, D(0) => 
                           NPC_Dec_0_port, Q(31) => NPC_ex_31_port, Q(30) => 
                           NPC_ex_30_port, Q(29) => NPC_ex_29_port, Q(28) => 
                           NPC_ex_28_port, Q(27) => NPC_ex_27_port, Q(26) => 
                           NPC_ex_26_port, Q(25) => NPC_ex_25_port, Q(24) => 
                           NPC_ex_24_port, Q(23) => NPC_ex_23_port, Q(22) => 
                           NPC_ex_22_port, Q(21) => NPC_ex_21_port, Q(20) => 
                           NPC_ex_20_port, Q(19) => NPC_ex_19_port, Q(18) => 
                           NPC_ex_18_port, Q(17) => NPC_ex_17_port, Q(16) => 
                           NPC_ex_16_port, Q(15) => NPC_ex_15_port, Q(14) => 
                           NPC_ex_14_port, Q(13) => NPC_ex_13_port, Q(12) => 
                           NPC_ex_12_port, Q(11) => NPC_ex_11_port, Q(10) => 
                           NPC_ex_10_port, Q(9) => NPC_ex_9_port, Q(8) => 
                           NPC_ex_8_port, Q(7) => NPC_ex_7_port, Q(6) => 
                           NPC_ex_6_port, Q(5) => NPC_ex_5_port, Q(4) => 
                           NPC_ex_4_port, Q(3) => NPC_ex_3_port, Q(2) => 
                           NPC_ex_2_port, Q(1) => NPC_ex_1_port, Q(0) => 
                           NPC_ex_0_port);
   pipeline_A2 : regFFD_NBIT32_9 port map( CK => CLK, RESET => n9, ENABLE => 
                           RF1, D(31) => regA_31_port, D(30) => regA_30_port, 
                           D(29) => regA_29_port, D(28) => regA_28_port, D(27) 
                           => regA_27_port, D(26) => regA_26_port, D(25) => 
                           regA_25_port, D(24) => regA_24_port, D(23) => 
                           regA_23_port, D(22) => regA_22_port, D(21) => 
                           regA_21_port, D(20) => regA_20_port, D(19) => 
                           regA_19_port, D(18) => regA_18_port, D(17) => 
                           regA_17_port, D(16) => regA_16_port, D(15) => 
                           regA_15_port, D(14) => regA_14_port, D(13) => 
                           regA_13_port, D(12) => regA_12_port, D(11) => 
                           regA_11_port, D(10) => regA_10_port, D(9) => 
                           regA_9_port, D(8) => regA_8_port, D(7) => 
                           regA_7_port, D(6) => regA_6_port, D(5) => 
                           regA_5_port, D(4) => regA_4_port, D(3) => 
                           regA_3_port, D(2) => regA_2_port, D(1) => 
                           regA_1_port, D(0) => regA_0_port, Q(31) => 
                           regA_ex_31_port, Q(30) => regA_ex_30_port, Q(29) => 
                           regA_ex_29_port, Q(28) => regA_ex_28_port, Q(27) => 
                           regA_ex_27_port, Q(26) => regA_ex_26_port, Q(25) => 
                           regA_ex_25_port, Q(24) => regA_ex_24_port, Q(23) => 
                           regA_ex_23_port, Q(22) => regA_ex_22_port, Q(21) => 
                           regA_ex_21_port, Q(20) => regA_ex_20_port, Q(19) => 
                           regA_ex_19_port, Q(18) => regA_ex_18_port, Q(17) => 
                           regA_ex_17_port, Q(16) => regA_ex_16_port, Q(15) => 
                           regA_ex_15_port, Q(14) => regA_ex_14_port, Q(13) => 
                           regA_ex_13_port, Q(12) => regA_ex_12_port, Q(11) => 
                           regA_ex_11_port, Q(10) => regA_ex_10_port, Q(9) => 
                           regA_ex_9_port, Q(8) => regA_ex_8_port, Q(7) => 
                           regA_ex_7_port, Q(6) => regA_ex_6_port, Q(5) => 
                           regA_ex_5_port, Q(4) => regA_ex_4_port, Q(3) => 
                           regA_ex_3_port, Q(2) => regA_ex_2_port, Q(1) => 
                           regA_ex_1_port, Q(0) => regA_ex_0_port);
   pipeline_B2 : regFFD_NBIT32_8 port map( CK => CLK, RESET => n9, ENABLE => 
                           RF2, D(31) => regB_31_port, D(30) => regB_30_port, 
                           D(29) => regB_29_port, D(28) => regB_28_port, D(27) 
                           => regB_27_port, D(26) => regB_26_port, D(25) => 
                           regB_25_port, D(24) => regB_24_port, D(23) => 
                           regB_23_port, D(22) => regB_22_port, D(21) => 
                           regB_21_port, D(20) => regB_20_port, D(19) => 
                           regB_19_port, D(18) => regB_18_port, D(17) => 
                           regB_17_port, D(16) => regB_16_port, D(15) => 
                           regB_15_port, D(14) => regB_14_port, D(13) => 
                           regB_13_port, D(12) => regB_12_port, D(11) => 
                           regB_11_port, D(10) => regB_10_port, D(9) => 
                           regB_9_port, D(8) => regB_8_port, D(7) => 
                           regB_7_port, D(6) => regB_6_port, D(5) => 
                           regB_5_port, D(4) => regB_4_port, D(3) => 
                           regB_3_port, D(2) => regB_2_port, D(1) => 
                           regB_1_port, D(0) => regB_0_port, Q(31) => 
                           regB_ex_31_port, Q(30) => regB_ex_30_port, Q(29) => 
                           regB_ex_29_port, Q(28) => regB_ex_28_port, Q(27) => 
                           regB_ex_27_port, Q(26) => regB_ex_26_port, Q(25) => 
                           regB_ex_25_port, Q(24) => regB_ex_24_port, Q(23) => 
                           regB_ex_23_port, Q(22) => regB_ex_22_port, Q(21) => 
                           regB_ex_21_port, Q(20) => regB_ex_20_port, Q(19) => 
                           regB_ex_19_port, Q(18) => regB_ex_18_port, Q(17) => 
                           regB_ex_17_port, Q(16) => regB_ex_16_port, Q(15) => 
                           regB_ex_15_port, Q(14) => regB_ex_14_port, Q(13) => 
                           regB_ex_13_port, Q(12) => regB_ex_12_port, Q(11) => 
                           regB_ex_11_port, Q(10) => regB_ex_10_port, Q(9) => 
                           regB_ex_9_port, Q(8) => regB_ex_8_port, Q(7) => 
                           regB_ex_7_port, Q(6) => regB_ex_6_port, Q(5) => 
                           regB_ex_5_port, Q(4) => regB_ex_4_port, Q(3) => 
                           regB_ex_3_port, Q(2) => regB_ex_2_port, Q(1) => 
                           regB_ex_1_port, Q(0) => regB_ex_0_port);
   pipeline_IMM2 : regFFD_NBIT32_7 port map( CK => CLK, RESET => n9, ENABLE => 
                           regImm_LATCH_EN, D(31) => Imm_31_port, D(30) => 
                           Imm_30_port, D(29) => Imm_29_port, D(28) => 
                           Imm_28_port, D(27) => Imm_27_port, D(26) => 
                           Imm_26_port, D(25) => Imm_25_port, D(24) => 
                           Imm_24_port, D(23) => Imm_23_port, D(22) => 
                           Imm_22_port, D(21) => Imm_21_port, D(20) => 
                           Imm_20_port, D(19) => Imm_19_port, D(18) => 
                           Imm_18_port, D(17) => Imm_17_port, D(16) => 
                           Imm_16_port, D(15) => Imm_15_port, D(14) => 
                           Imm_14_port, D(13) => Imm_13_port, D(12) => 
                           Imm_12_port, D(11) => Imm_11_port, D(10) => 
                           Imm_10_port, D(9) => Imm_9_port, D(8) => Imm_8_port,
                           D(7) => Imm_7_port, D(6) => Imm_6_port, D(5) => 
                           Imm_5_port, D(4) => Imm_4_port, D(3) => Imm_3_port, 
                           D(2) => Imm_2_port, D(1) => Imm_1_port, D(0) => 
                           Imm_0_port, Q(31) => Imm_ex_31_port, Q(30) => 
                           Imm_ex_30_port, Q(29) => Imm_ex_29_port, Q(28) => 
                           Imm_ex_28_port, Q(27) => Imm_ex_27_port, Q(26) => 
                           Imm_ex_26_port, Q(25) => Imm_ex_25_port, Q(24) => 
                           Imm_ex_24_port, Q(23) => Imm_ex_23_port, Q(22) => 
                           Imm_ex_22_port, Q(21) => Imm_ex_21_port, Q(20) => 
                           Imm_ex_20_port, Q(19) => Imm_ex_19_port, Q(18) => 
                           Imm_ex_18_port, Q(17) => Imm_ex_17_port, Q(16) => 
                           Imm_ex_16_port, Q(15) => Imm_ex_15_port, Q(14) => 
                           Imm_ex_14_port, Q(13) => Imm_ex_13_port, Q(12) => 
                           Imm_ex_12_port, Q(11) => Imm_ex_11_port, Q(10) => 
                           Imm_ex_10_port, Q(9) => Imm_ex_9_port, Q(8) => 
                           Imm_ex_8_port, Q(7) => Imm_ex_7_port, Q(6) => 
                           Imm_ex_6_port, Q(5) => Imm_ex_5_port, Q(4) => 
                           Imm_ex_4_port, Q(3) => Imm_ex_3_port, Q(2) => 
                           Imm_ex_2_port, Q(1) => Imm_ex_1_port, Q(0) => 
                           Imm_ex_0_port);
   pipeline_RD2 : regFFD_NBIT5_0 port map( CK => CLK, RESET => n8, ENABLE => 
                           X_Logic1_port, D(4) => RD_4_port, D(3) => RD_3_port,
                           D(2) => RD_2_port, D(1) => RD_1_port, D(0) => 
                           RD_0_port, Q(4) => RD_ex_4_port, Q(3) => 
                           RD_ex_3_port, Q(2) => RD_ex_2_port, Q(1) => 
                           RD_ex_1_port, Q(0) => RD_ex_0_port);
   pipeline_wr_signal : FF_7 port map( CLK => CLK, RESET => n9, EN => 
                           X_Logic1_port, D => n12, Q => wr_signal_exe);
   pipeline_IR2 : regFFD_NBIT6_0 port map( CK => CLK, RESET => n8, ENABLE => 
                           X_Logic1_port, D(5) => IR_Dec_31_port, D(4) => n1, 
                           D(3) => n2, D(2) => IR_Dec_28_port, D(1) => 
                           IR_Dec_27_port, D(0) => IR_Dec_26_port, Q(5) => 
                           IR_26_ex_5_port, Q(4) => IR_26_ex_4_port, Q(3) => 
                           IR_26_ex_3_port, Q(2) => IR_26_ex_2_port, Q(1) => 
                           IR_26_ex_1_port, Q(0) => IR_26_ex_0_port);
   pipeline_LHI2 : regFFD_NBIT32_6 port map( CK => CLK, RESET => n9, ENABLE => 
                           X_Logic1_port, D(31) => Imm_15_port, D(30) => 
                           Imm_14_port, D(29) => Imm_13_port, D(28) => 
                           Imm_12_port, D(27) => Imm_11_port, D(26) => 
                           Imm_10_port, D(25) => Imm_9_port, D(24) => 
                           Imm_8_port, D(23) => Imm_7_port, D(22) => Imm_6_port
                           , D(21) => Imm_5_port, D(20) => Imm_4_port, D(19) =>
                           Imm_3_port, D(18) => Imm_2_port, D(17) => Imm_1_port
                           , D(16) => Imm_0_port, D(15) => X_Logic0_port, D(14)
                           => X_Logic0_port, D(13) => X_Logic0_port, D(12) => 
                           X_Logic0_port, D(11) => X_Logic0_port, D(10) => 
                           X_Logic0_port, D(9) => X_Logic0_port, D(8) => 
                           X_Logic0_port, D(7) => X_Logic0_port, D(6) => 
                           X_Logic0_port, D(5) => X_Logic0_port, D(4) => 
                           X_Logic0_port, D(3) => X_Logic0_port, D(2) => 
                           X_Logic0_port, D(1) => X_Logic0_port, D(0) => 
                           X_Logic0_port, Q(31) => LHI_ex_31_port, Q(30) => 
                           LHI_ex_30_port, Q(29) => LHI_ex_29_port, Q(28) => 
                           LHI_ex_28_port, Q(27) => LHI_ex_27_port, Q(26) => 
                           LHI_ex_26_port, Q(25) => LHI_ex_25_port, Q(24) => 
                           LHI_ex_24_port, Q(23) => LHI_ex_23_port, Q(22) => 
                           LHI_ex_22_port, Q(21) => LHI_ex_21_port, Q(20) => 
                           LHI_ex_20_port, Q(19) => LHI_ex_19_port, Q(18) => 
                           LHI_ex_18_port, Q(17) => LHI_ex_17_port, Q(16) => 
                           LHI_ex_16_port, Q(15) => LHI_ex_15_port, Q(14) => 
                           LHI_ex_14_port, Q(13) => LHI_ex_13_port, Q(12) => 
                           LHI_ex_12_port, Q(11) => LHI_ex_11_port, Q(10) => 
                           LHI_ex_10_port, Q(9) => LHI_ex_9_port, Q(8) => 
                           LHI_ex_8_port, Q(7) => LHI_ex_7_port, Q(6) => 
                           LHI_ex_6_port, Q(5) => LHI_ex_5_port, Q(4) => 
                           LHI_ex_4_port, Q(3) => LHI_ex_3_port, Q(2) => 
                           LHI_ex_2_port, Q(1) => LHI_ex_1_port, Q(0) => 
                           LHI_ex_0_port);
   MUX_ALU_A : MUX21_GENERIC_NBIT32_6 port map( A(31) => NPC_ex_31_port, A(30) 
                           => NPC_ex_30_port, A(29) => NPC_ex_29_port, A(28) =>
                           NPC_ex_28_port, A(27) => NPC_ex_27_port, A(26) => 
                           NPC_ex_26_port, A(25) => NPC_ex_25_port, A(24) => 
                           NPC_ex_24_port, A(23) => NPC_ex_23_port, A(22) => 
                           NPC_ex_22_port, A(21) => NPC_ex_21_port, A(20) => 
                           NPC_ex_20_port, A(19) => NPC_ex_19_port, A(18) => 
                           NPC_ex_18_port, A(17) => NPC_ex_17_port, A(16) => 
                           NPC_ex_16_port, A(15) => NPC_ex_15_port, A(14) => 
                           NPC_ex_14_port, A(13) => NPC_ex_13_port, A(12) => 
                           NPC_ex_12_port, A(11) => NPC_ex_11_port, A(10) => 
                           NPC_ex_10_port, A(9) => NPC_ex_9_port, A(8) => 
                           NPC_ex_8_port, A(7) => NPC_ex_7_port, A(6) => 
                           NPC_ex_6_port, A(5) => NPC_ex_5_port, A(4) => 
                           NPC_ex_4_port, A(3) => NPC_ex_3_port, A(2) => 
                           NPC_ex_2_port, A(1) => NPC_ex_1_port, A(0) => 
                           NPC_ex_0_port, B(31) => regA_ex_31_port, B(30) => 
                           regA_ex_30_port, B(29) => regA_ex_29_port, B(28) => 
                           regA_ex_28_port, B(27) => regA_ex_27_port, B(26) => 
                           regA_ex_26_port, B(25) => regA_ex_25_port, B(24) => 
                           regA_ex_24_port, B(23) => regA_ex_23_port, B(22) => 
                           regA_ex_22_port, B(21) => regA_ex_21_port, B(20) => 
                           regA_ex_20_port, B(19) => regA_ex_19_port, B(18) => 
                           regA_ex_18_port, B(17) => regA_ex_17_port, B(16) => 
                           regA_ex_16_port, B(15) => regA_ex_15_port, B(14) => 
                           regA_ex_14_port, B(13) => regA_ex_13_port, B(12) => 
                           regA_ex_12_port, B(11) => regA_ex_11_port, B(10) => 
                           regA_ex_10_port, B(9) => regA_ex_9_port, B(8) => 
                           regA_ex_8_port, B(7) => regA_ex_7_port, B(6) => 
                           regA_ex_6_port, B(5) => regA_ex_5_port, B(4) => 
                           regA_ex_4_port, B(3) => regA_ex_3_port, B(2) => 
                           regA_ex_2_port, B(1) => regA_ex_1_port, B(0) => 
                           regA_ex_0_port, SEL => S1, Y(31) => 
                           input1_ALU_31_port, Y(30) => input1_ALU_30_port, 
                           Y(29) => input1_ALU_29_port, Y(28) => 
                           input1_ALU_28_port, Y(27) => input1_ALU_27_port, 
                           Y(26) => input1_ALU_26_port, Y(25) => 
                           input1_ALU_25_port, Y(24) => input1_ALU_24_port, 
                           Y(23) => input1_ALU_23_port, Y(22) => 
                           input1_ALU_22_port, Y(21) => input1_ALU_21_port, 
                           Y(20) => input1_ALU_20_port, Y(19) => 
                           input1_ALU_19_port, Y(18) => input1_ALU_18_port, 
                           Y(17) => input1_ALU_17_port, Y(16) => 
                           input1_ALU_16_port, Y(15) => input1_ALU_15_port, 
                           Y(14) => input1_ALU_14_port, Y(13) => 
                           input1_ALU_13_port, Y(12) => input1_ALU_12_port, 
                           Y(11) => input1_ALU_11_port, Y(10) => 
                           input1_ALU_10_port, Y(9) => input1_ALU_9_port, Y(8) 
                           => input1_ALU_8_port, Y(7) => input1_ALU_7_port, 
                           Y(6) => input1_ALU_6_port, Y(5) => input1_ALU_5_port
                           , Y(4) => input1_ALU_4_port, Y(3) => 
                           input1_ALU_3_port, Y(2) => input1_ALU_2_port, Y(1) 
                           => input1_ALU_1_port, Y(0) => input1_ALU_0_port);
   MUX_ALU_B : MUX21_GENERIC_NBIT32_5 port map( A(31) => Imm_ex_31_port, A(30) 
                           => Imm_ex_30_port, A(29) => Imm_ex_29_port, A(28) =>
                           Imm_ex_28_port, A(27) => Imm_ex_27_port, A(26) => 
                           Imm_ex_26_port, A(25) => Imm_ex_25_port, A(24) => 
                           Imm_ex_24_port, A(23) => Imm_ex_23_port, A(22) => 
                           Imm_ex_22_port, A(21) => Imm_ex_21_port, A(20) => 
                           Imm_ex_20_port, A(19) => Imm_ex_19_port, A(18) => 
                           Imm_ex_18_port, A(17) => Imm_ex_17_port, A(16) => 
                           Imm_ex_16_port, A(15) => Imm_ex_15_port, A(14) => 
                           Imm_ex_14_port, A(13) => Imm_ex_13_port, A(12) => 
                           Imm_ex_12_port, A(11) => Imm_ex_11_port, A(10) => 
                           Imm_ex_10_port, A(9) => Imm_ex_9_port, A(8) => 
                           Imm_ex_8_port, A(7) => Imm_ex_7_port, A(6) => 
                           Imm_ex_6_port, A(5) => Imm_ex_5_port, A(4) => 
                           Imm_ex_4_port, A(3) => Imm_ex_3_port, A(2) => 
                           Imm_ex_2_port, A(1) => Imm_ex_1_port, A(0) => 
                           Imm_ex_0_port, B(31) => regB_ex_31_port, B(30) => 
                           regB_ex_30_port, B(29) => regB_ex_29_port, B(28) => 
                           regB_ex_28_port, B(27) => regB_ex_27_port, B(26) => 
                           regB_ex_26_port, B(25) => regB_ex_25_port, B(24) => 
                           regB_ex_24_port, B(23) => regB_ex_23_port, B(22) => 
                           regB_ex_22_port, B(21) => regB_ex_21_port, B(20) => 
                           regB_ex_20_port, B(19) => regB_ex_19_port, B(18) => 
                           regB_ex_18_port, B(17) => regB_ex_17_port, B(16) => 
                           regB_ex_16_port, B(15) => regB_ex_15_port, B(14) => 
                           regB_ex_14_port, B(13) => regB_ex_13_port, B(12) => 
                           regB_ex_12_port, B(11) => regB_ex_11_port, B(10) => 
                           regB_ex_10_port, B(9) => regB_ex_9_port, B(8) => 
                           regB_ex_8_port, B(7) => regB_ex_7_port, B(6) => 
                           regB_ex_6_port, B(5) => regB_ex_5_port, B(4) => 
                           regB_ex_4_port, B(3) => regB_ex_3_port, B(2) => 
                           regB_ex_2_port, B(1) => regB_ex_1_port, B(0) => 
                           regB_ex_0_port, SEL => S2, Y(31) => 
                           input2_ALU_31_port, Y(30) => input2_ALU_30_port, 
                           Y(29) => input2_ALU_29_port, Y(28) => 
                           input2_ALU_28_port, Y(27) => input2_ALU_27_port, 
                           Y(26) => input2_ALU_26_port, Y(25) => 
                           input2_ALU_25_port, Y(24) => input2_ALU_24_port, 
                           Y(23) => input2_ALU_23_port, Y(22) => 
                           input2_ALU_22_port, Y(21) => input2_ALU_21_port, 
                           Y(20) => input2_ALU_20_port, Y(19) => 
                           input2_ALU_19_port, Y(18) => input2_ALU_18_port, 
                           Y(17) => input2_ALU_17_port, Y(16) => 
                           input2_ALU_16_port, Y(15) => input2_ALU_15_port, 
                           Y(14) => input2_ALU_14_port, Y(13) => 
                           input2_ALU_13_port, Y(12) => input2_ALU_12_port, 
                           Y(11) => input2_ALU_11_port, Y(10) => 
                           input2_ALU_10_port, Y(9) => input2_ALU_9_port, Y(8) 
                           => input2_ALU_8_port, Y(7) => input2_ALU_7_port, 
                           Y(6) => input2_ALU_6_port, Y(5) => input2_ALU_5_port
                           , Y(4) => input2_ALU_4_port, Y(3) => 
                           input2_ALU_3_port, Y(2) => input2_ALU_2_port, Y(1) 
                           => input2_ALU_1_port, Y(0) => input2_ALU_0_port);
   ALU_OP : ALU_N32 port map( CLK => CLK, FUNC(0) => instruction_alu(0), 
                           FUNC(1) => instruction_alu(1), FUNC(2) => 
                           instruction_alu(2), FUNC(3) => instruction_alu(3), 
                           FUNC(4) => instruction_alu(4), FUNC(5) => 
                           instruction_alu(5), DATA1(31) => input1_ALU_31_port,
                           DATA1(30) => input1_ALU_30_port, DATA1(29) => 
                           input1_ALU_29_port, DATA1(28) => input1_ALU_28_port,
                           DATA1(27) => input1_ALU_27_port, DATA1(26) => 
                           input1_ALU_26_port, DATA1(25) => input1_ALU_25_port,
                           DATA1(24) => input1_ALU_24_port, DATA1(23) => 
                           input1_ALU_23_port, DATA1(22) => input1_ALU_22_port,
                           DATA1(21) => input1_ALU_21_port, DATA1(20) => 
                           input1_ALU_20_port, DATA1(19) => input1_ALU_19_port,
                           DATA1(18) => input1_ALU_18_port, DATA1(17) => 
                           input1_ALU_17_port, DATA1(16) => input1_ALU_16_port,
                           DATA1(15) => input1_ALU_15_port, DATA1(14) => 
                           input1_ALU_14_port, DATA1(13) => input1_ALU_13_port,
                           DATA1(12) => input1_ALU_12_port, DATA1(11) => 
                           input1_ALU_11_port, DATA1(10) => input1_ALU_10_port,
                           DATA1(9) => input1_ALU_9_port, DATA1(8) => 
                           input1_ALU_8_port, DATA1(7) => input1_ALU_7_port, 
                           DATA1(6) => input1_ALU_6_port, DATA1(5) => 
                           input1_ALU_5_port, DATA1(4) => input1_ALU_4_port, 
                           DATA1(3) => input1_ALU_3_port, DATA1(2) => 
                           input1_ALU_2_port, DATA1(1) => input1_ALU_1_port, 
                           DATA1(0) => input1_ALU_0_port, DATA2(31) => 
                           input2_ALU_31_port, DATA2(30) => input2_ALU_30_port,
                           DATA2(29) => input2_ALU_29_port, DATA2(28) => 
                           input2_ALU_28_port, DATA2(27) => input2_ALU_27_port,
                           DATA2(26) => input2_ALU_26_port, DATA2(25) => 
                           input2_ALU_25_port, DATA2(24) => input2_ALU_24_port,
                           DATA2(23) => input2_ALU_23_port, DATA2(22) => 
                           input2_ALU_22_port, DATA2(21) => input2_ALU_21_port,
                           DATA2(20) => input2_ALU_20_port, DATA2(19) => 
                           input2_ALU_19_port, DATA2(18) => input2_ALU_18_port,
                           DATA2(17) => input2_ALU_17_port, DATA2(16) => 
                           input2_ALU_16_port, DATA2(15) => input2_ALU_15_port,
                           DATA2(14) => input2_ALU_14_port, DATA2(13) => 
                           input2_ALU_13_port, DATA2(12) => input2_ALU_12_port,
                           DATA2(11) => input2_ALU_11_port, DATA2(10) => 
                           input2_ALU_10_port, DATA2(9) => input2_ALU_9_port, 
                           DATA2(8) => input2_ALU_8_port, DATA2(7) => 
                           input2_ALU_7_port, DATA2(6) => input2_ALU_6_port, 
                           DATA2(5) => input2_ALU_5_port, DATA2(4) => 
                           input2_ALU_4_port, DATA2(3) => input2_ALU_3_port, 
                           DATA2(2) => input2_ALU_2_port, DATA2(1) => 
                           input2_ALU_1_port, DATA2(0) => input2_ALU_0_port, 
                           OUT_ALU(31) => ALU_out_31_port, OUT_ALU(30) => 
                           ALU_out_30_port, OUT_ALU(29) => ALU_out_29_port, 
                           OUT_ALU(28) => ALU_out_28_port, OUT_ALU(27) => 
                           ALU_out_27_port, OUT_ALU(26) => ALU_out_26_port, 
                           OUT_ALU(25) => ALU_out_25_port, OUT_ALU(24) => 
                           ALU_out_24_port, OUT_ALU(23) => ALU_out_23_port, 
                           OUT_ALU(22) => ALU_out_22_port, OUT_ALU(21) => 
                           ALU_out_21_port, OUT_ALU(20) => ALU_out_20_port, 
                           OUT_ALU(19) => ALU_out_19_port, OUT_ALU(18) => 
                           ALU_out_18_port, OUT_ALU(17) => ALU_out_17_port, 
                           OUT_ALU(16) => ALU_out_16_port, OUT_ALU(15) => 
                           ALU_out_15_port, OUT_ALU(14) => ALU_out_14_port, 
                           OUT_ALU(13) => ALU_out_13_port, OUT_ALU(12) => 
                           ALU_out_12_port, OUT_ALU(11) => ALU_out_11_port, 
                           OUT_ALU(10) => ALU_out_10_port, OUT_ALU(9) => 
                           ALU_out_9_port, OUT_ALU(8) => ALU_out_8_port, 
                           OUT_ALU(7) => ALU_out_7_port, OUT_ALU(6) => 
                           ALU_out_6_port, OUT_ALU(5) => ALU_out_5_port, 
                           OUT_ALU(4) => ALU_out_4_port, OUT_ALU(3) => 
                           ALU_out_3_port, OUT_ALU(2) => ALU_out_2_port, 
                           OUT_ALU(1) => ALU_out_1_port, OUT_ALU(0) => 
                           ALU_out_0_port);
   ZERO_OP : zero_eval_NBIT32 port map( input(31) => regA_ex_31_port, input(30)
                           => regA_ex_30_port, input(29) => regA_ex_29_port, 
                           input(28) => regA_ex_28_port, input(27) => 
                           regA_ex_27_port, input(26) => regA_ex_26_port, 
                           input(25) => regA_ex_25_port, input(24) => 
                           regA_ex_24_port, input(23) => regA_ex_23_port, 
                           input(22) => regA_ex_22_port, input(21) => 
                           regA_ex_21_port, input(20) => regA_ex_20_port, 
                           input(19) => regA_ex_19_port, input(18) => 
                           regA_ex_18_port, input(17) => regA_ex_17_port, 
                           input(16) => regA_ex_16_port, input(15) => 
                           regA_ex_15_port, input(14) => regA_ex_14_port, 
                           input(13) => regA_ex_13_port, input(12) => 
                           regA_ex_12_port, input(11) => regA_ex_11_port, 
                           input(10) => regA_ex_10_port, input(9) => 
                           regA_ex_9_port, input(8) => regA_ex_8_port, input(7)
                           => regA_ex_7_port, input(6) => regA_ex_6_port, 
                           input(5) => regA_ex_5_port, input(4) => 
                           regA_ex_4_port, input(3) => regA_ex_3_port, input(2)
                           => regA_ex_2_port, input(1) => regA_ex_1_port, 
                           input(0) => regA_ex_0_port, res => is_zero);
   COND_OP : COND_BT_NBIT32 port map( ZERO_BIT => is_zero, OPCODE_0 => 
                           IR_26_ex_0_port, branch_op => branch_cond, con_sign 
                           => cond);
   MUX_alu_out : MUX21_GENERIC_NBIT32_4 port map( A(31) => LHI_ex_31_port, 
                           A(30) => LHI_ex_30_port, A(29) => LHI_ex_29_port, 
                           A(28) => LHI_ex_28_port, A(27) => LHI_ex_27_port, 
                           A(26) => LHI_ex_26_port, A(25) => LHI_ex_25_port, 
                           A(24) => LHI_ex_24_port, A(23) => LHI_ex_23_port, 
                           A(22) => LHI_ex_22_port, A(21) => LHI_ex_21_port, 
                           A(20) => LHI_ex_20_port, A(19) => LHI_ex_19_port, 
                           A(18) => LHI_ex_18_port, A(17) => LHI_ex_17_port, 
                           A(16) => LHI_ex_16_port, A(15) => LHI_ex_15_port, 
                           A(14) => LHI_ex_14_port, A(13) => LHI_ex_13_port, 
                           A(12) => LHI_ex_12_port, A(11) => LHI_ex_11_port, 
                           A(10) => LHI_ex_10_port, A(9) => LHI_ex_9_port, A(8)
                           => LHI_ex_8_port, A(7) => LHI_ex_7_port, A(6) => 
                           LHI_ex_6_port, A(5) => LHI_ex_5_port, A(4) => 
                           LHI_ex_4_port, A(3) => LHI_ex_3_port, A(2) => 
                           LHI_ex_2_port, A(1) => LHI_ex_1_port, A(0) => 
                           LHI_ex_0_port, B(31) => ALU_out_31_port, B(30) => 
                           ALU_out_30_port, B(29) => ALU_out_29_port, B(28) => 
                           ALU_out_28_port, B(27) => ALU_out_27_port, B(26) => 
                           ALU_out_26_port, B(25) => ALU_out_25_port, B(24) => 
                           ALU_out_24_port, B(23) => ALU_out_23_port, B(22) => 
                           ALU_out_22_port, B(21) => ALU_out_21_port, B(20) => 
                           ALU_out_20_port, B(19) => ALU_out_19_port, B(18) => 
                           ALU_out_18_port, B(17) => ALU_out_17_port, B(16) => 
                           ALU_out_16_port, B(15) => ALU_out_15_port, B(14) => 
                           ALU_out_14_port, B(13) => ALU_out_13_port, B(12) => 
                           ALU_out_12_port, B(11) => ALU_out_11_port, B(10) => 
                           ALU_out_10_port, B(9) => ALU_out_9_port, B(8) => 
                           ALU_out_8_port, B(7) => ALU_out_7_port, B(6) => 
                           ALU_out_6_port, B(5) => ALU_out_5_port, B(4) => 
                           ALU_out_4_port, B(3) => ALU_out_3_port, B(2) => 
                           ALU_out_2_port, B(1) => ALU_out_1_port, B(0) => 
                           ALU_out_0_port, SEL => lhi_sel, Y(31) => 
                           ALU_ex_31_port, Y(30) => ALU_ex_30_port, Y(29) => 
                           ALU_ex_29_port, Y(28) => ALU_ex_28_port, Y(27) => 
                           ALU_ex_27_port, Y(26) => ALU_ex_26_port, Y(25) => 
                           ALU_ex_25_port, Y(24) => ALU_ex_24_port, Y(23) => 
                           ALU_ex_23_port, Y(22) => ALU_ex_22_port, Y(21) => 
                           ALU_ex_21_port, Y(20) => ALU_ex_20_port, Y(19) => 
                           ALU_ex_19_port, Y(18) => ALU_ex_18_port, Y(17) => 
                           ALU_ex_17_port, Y(16) => ALU_ex_16_port, Y(15) => 
                           ALU_ex_15_port, Y(14) => ALU_ex_14_port, Y(13) => 
                           ALU_ex_13_port, Y(12) => ALU_ex_12_port, Y(11) => 
                           ALU_ex_11_port, Y(10) => ALU_ex_10_port, Y(9) => 
                           ALU_ex_9_port, Y(8) => ALU_ex_8_port, Y(7) => 
                           ALU_ex_7_port, Y(6) => ALU_ex_6_port, Y(5) => 
                           ALU_ex_5_port, Y(4) => ALU_ex_4_port, Y(3) => 
                           ALU_ex_3_port, Y(2) => ALU_ex_2_port, Y(1) => 
                           ALU_ex_1_port, Y(0) => ALU_ex_0_port);
   pipeline_sign3 : FF_6 port map( CLK => CLK, RESET => n9, EN => X_Logic1_port
                           , D => signed_op_ex, Q => signed_op_mem);
   pipeline_newpc3 : regFFD_NBIT32_5 port map( CK => CLK, RESET => n9, ENABLE 
                           => X_Logic1_port, D(31) => NPC_ex_31_port, D(30) => 
                           NPC_ex_30_port, D(29) => NPC_ex_29_port, D(28) => 
                           NPC_ex_28_port, D(27) => NPC_ex_27_port, D(26) => 
                           NPC_ex_26_port, D(25) => NPC_ex_25_port, D(24) => 
                           NPC_ex_24_port, D(23) => NPC_ex_23_port, D(22) => 
                           NPC_ex_22_port, D(21) => NPC_ex_21_port, D(20) => 
                           NPC_ex_20_port, D(19) => NPC_ex_19_port, D(18) => 
                           NPC_ex_18_port, D(17) => NPC_ex_17_port, D(16) => 
                           NPC_ex_16_port, D(15) => NPC_ex_15_port, D(14) => 
                           NPC_ex_14_port, D(13) => NPC_ex_13_port, D(12) => 
                           NPC_ex_12_port, D(11) => NPC_ex_11_port, D(10) => 
                           NPC_ex_10_port, D(9) => NPC_ex_9_port, D(8) => 
                           NPC_ex_8_port, D(7) => NPC_ex_7_port, D(6) => 
                           NPC_ex_6_port, D(5) => NPC_ex_5_port, D(4) => 
                           NPC_ex_4_port, D(3) => NPC_ex_3_port, D(2) => 
                           NPC_ex_2_port, D(1) => NPC_ex_1_port, D(0) => 
                           NPC_ex_0_port, Q(31) => NPC_mem_31_port, Q(30) => 
                           NPC_mem_30_port, Q(29) => NPC_mem_29_port, Q(28) => 
                           NPC_mem_28_port, Q(27) => NPC_mem_27_port, Q(26) => 
                           NPC_mem_26_port, Q(25) => NPC_mem_25_port, Q(24) => 
                           NPC_mem_24_port, Q(23) => NPC_mem_23_port, Q(22) => 
                           NPC_mem_22_port, Q(21) => NPC_mem_21_port, Q(20) => 
                           NPC_mem_20_port, Q(19) => NPC_mem_19_port, Q(18) => 
                           NPC_mem_18_port, Q(17) => NPC_mem_17_port, Q(16) => 
                           NPC_mem_16_port, Q(15) => NPC_mem_15_port, Q(14) => 
                           NPC_mem_14_port, Q(13) => NPC_mem_13_port, Q(12) => 
                           NPC_mem_12_port, Q(11) => NPC_mem_11_port, Q(10) => 
                           NPC_mem_10_port, Q(9) => NPC_mem_9_port, Q(8) => 
                           NPC_mem_8_port, Q(7) => NPC_mem_7_port, Q(6) => 
                           NPC_mem_6_port, Q(5) => NPC_mem_5_port, Q(4) => 
                           NPC_mem_4_port, Q(3) => NPC_mem_3_port, Q(2) => 
                           NPC_mem_2_port, Q(1) => NPC_mem_1_port, Q(0) => 
                           NPC_mem_0_port);
   pipeline_cond3 : FF_5 port map( CLK => CLK, RESET => n9, EN => X_Logic1_port
                           , D => cond, Q => cond_mem);
   pipeline_B3 : regFFD_NBIT32_4 port map( CK => CLK, RESET => n8, ENABLE => 
                           X_Logic1_port, D(31) => regB_ex_31_port, D(30) => 
                           regB_ex_30_port, D(29) => regB_ex_29_port, D(28) => 
                           regB_ex_28_port, D(27) => regB_ex_27_port, D(26) => 
                           regB_ex_26_port, D(25) => regB_ex_25_port, D(24) => 
                           regB_ex_24_port, D(23) => regB_ex_23_port, D(22) => 
                           regB_ex_22_port, D(21) => regB_ex_21_port, D(20) => 
                           regB_ex_20_port, D(19) => regB_ex_19_port, D(18) => 
                           regB_ex_18_port, D(17) => regB_ex_17_port, D(16) => 
                           regB_ex_16_port, D(15) => regB_ex_15_port, D(14) => 
                           regB_ex_14_port, D(13) => regB_ex_13_port, D(12) => 
                           regB_ex_12_port, D(11) => regB_ex_11_port, D(10) => 
                           regB_ex_10_port, D(9) => regB_ex_9_port, D(8) => 
                           regB_ex_8_port, D(7) => regB_ex_7_port, D(6) => 
                           regB_ex_6_port, D(5) => regB_ex_5_port, D(4) => 
                           regB_ex_4_port, D(3) => regB_ex_3_port, D(2) => 
                           regB_ex_2_port, D(1) => regB_ex_1_port, D(0) => 
                           regB_ex_0_port, Q(31) => regB_mem_31_port, Q(30) => 
                           regB_mem_30_port, Q(29) => regB_mem_29_port, Q(28) 
                           => regB_mem_28_port, Q(27) => regB_mem_27_port, 
                           Q(26) => regB_mem_26_port, Q(25) => regB_mem_25_port
                           , Q(24) => regB_mem_24_port, Q(23) => 
                           regB_mem_23_port, Q(22) => regB_mem_22_port, Q(21) 
                           => regB_mem_21_port, Q(20) => regB_mem_20_port, 
                           Q(19) => regB_mem_19_port, Q(18) => regB_mem_18_port
                           , Q(17) => regB_mem_17_port, Q(16) => 
                           regB_mem_16_port, Q(15) => regB_mem_15_port, Q(14) 
                           => regB_mem_14_port, Q(13) => regB_mem_13_port, 
                           Q(12) => regB_mem_12_port, Q(11) => regB_mem_11_port
                           , Q(10) => regB_mem_10_port, Q(9) => regB_mem_9_port
                           , Q(8) => regB_mem_8_port, Q(7) => regB_mem_7_port, 
                           Q(6) => regB_mem_6_port, Q(5) => regB_mem_5_port, 
                           Q(4) => regB_mem_4_port, Q(3) => regB_mem_3_port, 
                           Q(2) => regB_mem_2_port, Q(1) => regB_mem_1_port, 
                           Q(0) => regB_mem_0_port);
   pipeline_RD3 : regFFD_NBIT5_2 port map( CK => CLK, RESET => n8, ENABLE => 
                           X_Logic1_port, D(4) => RD_ex_4_port, D(3) => 
                           RD_ex_3_port, D(2) => RD_ex_2_port, D(1) => 
                           RD_ex_1_port, D(0) => RD_ex_0_port, Q(4) => 
                           RD_mem_4_port, Q(3) => RD_mem_3_port, Q(2) => 
                           RD_mem_2_port, Q(1) => RD_mem_1_port, Q(0) => 
                           RD_mem_0_port);
   pipeline_wr_signal2 : FF_4 port map( CLK => CLK, RESET => n9, EN => 
                           X_Logic1_port, D => wr_signal_exe, Q => 
                           wr_signal_mem);
   pipeline_IR3 : regFFD_NBIT6_1 port map( CK => CLK, RESET => n8, ENABLE => 
                           X_Logic1_port, D(5) => IR_26_ex_5_port, D(4) => 
                           IR_26_ex_4_port, D(3) => IR_26_ex_3_port, D(2) => 
                           IR_26_ex_2_port, D(1) => IR_26_ex_1_port, D(0) => 
                           IR_26_ex_0_port, Q(5) => IR_26_mem_5_port, Q(4) => 
                           IR_26_mem_4_port, Q(3) => IR_26_mem_3_port, Q(2) => 
                           IR_26_mem_2_port, Q(1) => IR_26_mem_1_port, Q(0) => 
                           IR_26_mem_0_port);
   MUX_PC : MUX21_GENERIC_NBIT32_3 port map( A(31) => ALU_ex_31_port, A(30) => 
                           ALU_ex_30_port, A(29) => ALU_ex_29_port, A(28) => 
                           ALU_ex_28_port, A(27) => ALU_ex_27_port, A(26) => 
                           ALU_ex_26_port, A(25) => ALU_ex_25_port, A(24) => 
                           ALU_ex_24_port, A(23) => ALU_ex_23_port, A(22) => 
                           ALU_ex_22_port, A(21) => ALU_ex_21_port, A(20) => 
                           ALU_ex_20_port, A(19) => ALU_ex_19_port, A(18) => 
                           ALU_ex_18_port, A(17) => ALU_ex_17_port, A(16) => 
                           ALU_ex_16_port, A(15) => ALU_ex_15_port, A(14) => 
                           ALU_ex_14_port, A(13) => ALU_ex_13_port, A(12) => 
                           ALU_ex_12_port, A(11) => ALU_ex_11_port, A(10) => 
                           ALU_ex_10_port, A(9) => ALU_ex_9_port, A(8) => 
                           ALU_ex_8_port, A(7) => ALU_ex_7_port, A(6) => 
                           ALU_ex_6_port, A(5) => ALU_ex_5_port, A(4) => 
                           ALU_ex_4_port, A(3) => ALU_ex_3_port, A(2) => 
                           ALU_ex_2_port, A(1) => ALU_ex_1_port, A(0) => 
                           ALU_ex_0_port, B(31) => NPC_mem_31_port, B(30) => 
                           NPC_mem_30_port, B(29) => NPC_mem_29_port, B(28) => 
                           NPC_mem_28_port, B(27) => NPC_mem_27_port, B(26) => 
                           NPC_mem_26_port, B(25) => NPC_mem_25_port, B(24) => 
                           NPC_mem_24_port, B(23) => NPC_mem_23_port, B(22) => 
                           NPC_mem_22_port, B(21) => NPC_mem_21_port, B(20) => 
                           NPC_mem_20_port, B(19) => NPC_mem_19_port, B(18) => 
                           NPC_mem_18_port, B(17) => NPC_mem_17_port, B(16) => 
                           NPC_mem_16_port, B(15) => NPC_mem_15_port, B(14) => 
                           NPC_mem_14_port, B(13) => NPC_mem_13_port, B(12) => 
                           NPC_mem_12_port, B(11) => NPC_mem_11_port, B(10) => 
                           NPC_mem_10_port, B(9) => NPC_mem_9_port, B(8) => 
                           NPC_mem_8_port, B(7) => NPC_mem_7_port, B(6) => 
                           NPC_mem_6_port, B(5) => NPC_mem_5_port, B(4) => 
                           NPC_mem_4_port, B(3) => NPC_mem_3_port, B(2) => 
                           NPC_mem_2_port, B(1) => NPC_mem_1_port, B(0) => 
                           NPC_mem_0_port, SEL => sel_npc, Y(31) => 
                           PC_OUT_i_31_port, Y(30) => PC_OUT_i_30_port, Y(29) 
                           => PC_OUT_i_29_port, Y(28) => PC_OUT_i_28_port, 
                           Y(27) => PC_OUT_i_27_port, Y(26) => PC_OUT_i_26_port
                           , Y(25) => PC_OUT_i_25_port, Y(24) => 
                           PC_OUT_i_24_port, Y(23) => PC_OUT_i_23_port, Y(22) 
                           => PC_OUT_i_22_port, Y(21) => PC_OUT_i_21_port, 
                           Y(20) => PC_OUT_i_20_port, Y(19) => PC_OUT_i_19_port
                           , Y(18) => PC_OUT_i_18_port, Y(17) => 
                           PC_OUT_i_17_port, Y(16) => PC_OUT_i_16_port, Y(15) 
                           => PC_OUT_i_15_port, Y(14) => PC_OUT_i_14_port, 
                           Y(13) => PC_OUT_i_13_port, Y(12) => PC_OUT_i_12_port
                           , Y(11) => PC_OUT_i_11_port, Y(10) => 
                           PC_OUT_i_10_port, Y(9) => PC_OUT_i_9_port, Y(8) => 
                           PC_OUT_i_8_port, Y(7) => PC_OUT_i_7_port, Y(6) => 
                           PC_OUT_i_6_port, Y(5) => PC_OUT_i_5_port, Y(4) => 
                           PC_OUT_i_4_port, Y(3) => PC_OUT_i_3_port, Y(2) => 
                           PC_OUT_i_2_port, Y(1) => PC_OUT_i_1_port, Y(0) => 
                           PC_OUT_i_0_port);
   LOAD_DATA_OUT : load_data port map( data_in(31) => DATA_MEM_OUT(31), 
                           data_in(30) => DATA_MEM_OUT(30), data_in(29) => 
                           DATA_MEM_OUT(29), data_in(28) => DATA_MEM_OUT(28), 
                           data_in(27) => DATA_MEM_OUT(27), data_in(26) => 
                           DATA_MEM_OUT(26), data_in(25) => DATA_MEM_OUT(25), 
                           data_in(24) => DATA_MEM_OUT(24), data_in(23) => 
                           DATA_MEM_OUT(23), data_in(22) => DATA_MEM_OUT(22), 
                           data_in(21) => DATA_MEM_OUT(21), data_in(20) => 
                           DATA_MEM_OUT(20), data_in(19) => DATA_MEM_OUT(19), 
                           data_in(18) => DATA_MEM_OUT(18), data_in(17) => 
                           DATA_MEM_OUT(17), data_in(16) => DATA_MEM_OUT(16), 
                           data_in(15) => DATA_MEM_OUT(15), data_in(14) => 
                           DATA_MEM_OUT(14), data_in(13) => DATA_MEM_OUT(13), 
                           data_in(12) => DATA_MEM_OUT(12), data_in(11) => 
                           DATA_MEM_OUT(11), data_in(10) => DATA_MEM_OUT(10), 
                           data_in(9) => DATA_MEM_OUT(9), data_in(8) => 
                           DATA_MEM_OUT(8), data_in(7) => DATA_MEM_OUT(7), 
                           data_in(6) => DATA_MEM_OUT(6), data_in(5) => 
                           DATA_MEM_OUT(5), data_in(4) => DATA_MEM_OUT(4), 
                           data_in(3) => DATA_MEM_OUT(3), data_in(2) => 
                           DATA_MEM_OUT(2), data_in(1) => DATA_MEM_OUT(1), 
                           data_in(0) => DATA_MEM_OUT(0), signed_val => 
                           signed_op_mem, load_op => RM, load_type(1) => 
                           IR_26_mem_1_port, load_type(0) => IR_26_mem_0_port, 
                           data_out(31) => LMD_out_31_port, data_out(30) => 
                           LMD_out_30_port, data_out(29) => LMD_out_29_port, 
                           data_out(28) => LMD_out_28_port, data_out(27) => 
                           LMD_out_27_port, data_out(26) => LMD_out_26_port, 
                           data_out(25) => LMD_out_25_port, data_out(24) => 
                           LMD_out_24_port, data_out(23) => LMD_out_23_port, 
                           data_out(22) => LMD_out_22_port, data_out(21) => 
                           LMD_out_21_port, data_out(20) => LMD_out_20_port, 
                           data_out(19) => LMD_out_19_port, data_out(18) => 
                           LMD_out_18_port, data_out(17) => LMD_out_17_port, 
                           data_out(16) => LMD_out_16_port, data_out(15) => 
                           LMD_out_15_port, data_out(14) => LMD_out_14_port, 
                           data_out(13) => LMD_out_13_port, data_out(12) => 
                           LMD_out_12_port, data_out(11) => LMD_out_11_port, 
                           data_out(10) => LMD_out_10_port, data_out(9) => 
                           LMD_out_9_port, data_out(8) => LMD_out_8_port, 
                           data_out(7) => LMD_out_7_port, data_out(6) => 
                           LMD_out_6_port, data_out(5) => LMD_out_5_port, 
                           data_out(4) => LMD_out_4_port, data_out(3) => 
                           LMD_out_3_port, data_out(2) => LMD_out_2_port, 
                           data_out(1) => LMD_out_1_port, data_out(0) => 
                           LMD_out_0_port);
   pipeline_alu4 : regFFD_NBIT32_3 port map( CK => CLK, RESET => n8, ENABLE => 
                           X_Logic1_port, D(31) => ALU_ex_31_port, D(30) => 
                           ALU_ex_30_port, D(29) => ALU_ex_29_port, D(28) => 
                           ALU_ex_28_port, D(27) => ALU_ex_27_port, D(26) => 
                           ALU_ex_26_port, D(25) => ALU_ex_25_port, D(24) => 
                           ALU_ex_24_port, D(23) => ALU_ex_23_port, D(22) => 
                           ALU_ex_22_port, D(21) => ALU_ex_21_port, D(20) => 
                           ALU_ex_20_port, D(19) => ALU_ex_19_port, D(18) => 
                           ALU_ex_18_port, D(17) => ALU_ex_17_port, D(16) => 
                           ALU_ex_16_port, D(15) => ALU_ex_15_port, D(14) => 
                           ALU_ex_14_port, D(13) => ALU_ex_13_port, D(12) => 
                           ALU_ex_12_port, D(11) => ALU_ex_11_port, D(10) => 
                           ALU_ex_10_port, D(9) => ALU_ex_9_port, D(8) => 
                           ALU_ex_8_port, D(7) => ALU_ex_7_port, D(6) => 
                           ALU_ex_6_port, D(5) => ALU_ex_5_port, D(4) => 
                           ALU_ex_4_port, D(3) => ALU_ex_3_port, D(2) => 
                           ALU_ex_2_port, D(1) => ALU_ex_1_port, D(0) => 
                           ALU_ex_0_port, Q(31) => ALU_wb_31_port, Q(30) => 
                           ALU_wb_30_port, Q(29) => ALU_wb_29_port, Q(28) => 
                           ALU_wb_28_port, Q(27) => ALU_wb_27_port, Q(26) => 
                           ALU_wb_26_port, Q(25) => ALU_wb_25_port, Q(24) => 
                           ALU_wb_24_port, Q(23) => ALU_wb_23_port, Q(22) => 
                           ALU_wb_22_port, Q(21) => ALU_wb_21_port, Q(20) => 
                           ALU_wb_20_port, Q(19) => ALU_wb_19_port, Q(18) => 
                           ALU_wb_18_port, Q(17) => ALU_wb_17_port, Q(16) => 
                           ALU_wb_16_port, Q(15) => ALU_wb_15_port, Q(14) => 
                           ALU_wb_14_port, Q(13) => ALU_wb_13_port, Q(12) => 
                           ALU_wb_12_port, Q(11) => ALU_wb_11_port, Q(10) => 
                           ALU_wb_10_port, Q(9) => ALU_wb_9_port, Q(8) => 
                           ALU_wb_8_port, Q(7) => ALU_wb_7_port, Q(6) => 
                           ALU_wb_6_port, Q(5) => ALU_wb_5_port, Q(4) => 
                           ALU_wb_4_port, Q(3) => ALU_wb_3_port, Q(2) => 
                           ALU_wb_2_port, Q(1) => ALU_wb_1_port, Q(0) => 
                           ALU_wb_0_port);
   pipeline_LMD4 : regFFD_NBIT32_2 port map( CK => CLK, RESET => n8, ENABLE => 
                           RM, D(31) => LMD_out_31_port, D(30) => 
                           LMD_out_30_port, D(29) => LMD_out_29_port, D(28) => 
                           LMD_out_28_port, D(27) => LMD_out_27_port, D(26) => 
                           LMD_out_26_port, D(25) => LMD_out_25_port, D(24) => 
                           LMD_out_24_port, D(23) => LMD_out_23_port, D(22) => 
                           LMD_out_22_port, D(21) => LMD_out_21_port, D(20) => 
                           LMD_out_20_port, D(19) => LMD_out_19_port, D(18) => 
                           LMD_out_18_port, D(17) => LMD_out_17_port, D(16) => 
                           LMD_out_16_port, D(15) => LMD_out_15_port, D(14) => 
                           LMD_out_14_port, D(13) => LMD_out_13_port, D(12) => 
                           LMD_out_12_port, D(11) => LMD_out_11_port, D(10) => 
                           LMD_out_10_port, D(9) => LMD_out_9_port, D(8) => 
                           LMD_out_8_port, D(7) => LMD_out_7_port, D(6) => 
                           LMD_out_6_port, D(5) => LMD_out_5_port, D(4) => 
                           LMD_out_4_port, D(3) => LMD_out_3_port, D(2) => 
                           LMD_out_2_port, D(1) => LMD_out_1_port, D(0) => 
                           LMD_out_0_port, Q(31) => LMD_wb_31_port, Q(30) => 
                           LMD_wb_30_port, Q(29) => LMD_wb_29_port, Q(28) => 
                           LMD_wb_28_port, Q(27) => LMD_wb_27_port, Q(26) => 
                           LMD_wb_26_port, Q(25) => LMD_wb_25_port, Q(24) => 
                           LMD_wb_24_port, Q(23) => LMD_wb_23_port, Q(22) => 
                           LMD_wb_22_port, Q(21) => LMD_wb_21_port, Q(20) => 
                           LMD_wb_20_port, Q(19) => LMD_wb_19_port, Q(18) => 
                           LMD_wb_18_port, Q(17) => LMD_wb_17_port, Q(16) => 
                           LMD_wb_16_port, Q(15) => LMD_wb_15_port, Q(14) => 
                           LMD_wb_14_port, Q(13) => LMD_wb_13_port, Q(12) => 
                           LMD_wb_12_port, Q(11) => LMD_wb_11_port, Q(10) => 
                           LMD_wb_10_port, Q(9) => LMD_wb_9_port, Q(8) => 
                           LMD_wb_8_port, Q(7) => LMD_wb_7_port, Q(6) => 
                           LMD_wb_6_port, Q(5) => LMD_wb_5_port, Q(4) => 
                           LMD_wb_4_port, Q(3) => LMD_wb_3_port, Q(2) => 
                           LMD_wb_2_port, Q(1) => LMD_wb_1_port, Q(0) => 
                           LMD_wb_0_port);
   pipeline_RD4 : regFFD_NBIT5_1 port map( CK => CLK, RESET => n8, ENABLE => 
                           X_Logic1_port, D(4) => RD_mem_4_port, D(3) => 
                           RD_mem_3_port, D(2) => RD_mem_2_port, D(1) => 
                           RD_mem_1_port, D(0) => RD_mem_0_port, Q(4) => 
                           RD_wb_4_port, Q(3) => RD_wb_3_port, Q(2) => 
                           RD_wb_2_port, Q(1) => RD_wb_1_port, Q(0) => 
                           RD_wb_0_port);
   pipeline_wr_signal3 : FF_3 port map( CLK => CLK, RESET => n9, EN => 
                           X_Logic1_port, D => wr_signal_mem1, Q => 
                           wr_signal_wb);
   pipeline_WM : FF_2 port map( CLK => CLK, RESET => n9, EN => X_Logic1_port, D
                           => WM, Q => n_2357);
   pipeline_JAL : FF_1 port map( CLK => CLK, RESET => n9, EN => X_Logic1_port, 
                           D => sel_saved_reg, Q => sel_saved_reg_wb);
   pipeline_NPC_wb : regFFD_NBIT32_1 port map( CK => CLK, RESET => n8, ENABLE 
                           => X_Logic1_port, D(31) => NPC_mem_31_port, D(30) =>
                           NPC_mem_30_port, D(29) => NPC_mem_29_port, D(28) => 
                           NPC_mem_28_port, D(27) => NPC_mem_27_port, D(26) => 
                           NPC_mem_26_port, D(25) => NPC_mem_25_port, D(24) => 
                           NPC_mem_24_port, D(23) => NPC_mem_23_port, D(22) => 
                           NPC_mem_22_port, D(21) => NPC_mem_21_port, D(20) => 
                           NPC_mem_20_port, D(19) => NPC_mem_19_port, D(18) => 
                           NPC_mem_18_port, D(17) => NPC_mem_17_port, D(16) => 
                           NPC_mem_16_port, D(15) => NPC_mem_15_port, D(14) => 
                           NPC_mem_14_port, D(13) => NPC_mem_13_port, D(12) => 
                           NPC_mem_12_port, D(11) => NPC_mem_11_port, D(10) => 
                           NPC_mem_10_port, D(9) => NPC_mem_9_port, D(8) => 
                           NPC_mem_8_port, D(7) => NPC_mem_7_port, D(6) => 
                           NPC_mem_6_port, D(5) => NPC_mem_5_port, D(4) => 
                           NPC_mem_4_port, D(3) => NPC_mem_3_port, D(2) => 
                           NPC_mem_2_port, D(1) => NPC_mem_1_port, D(0) => 
                           NPC_mem_0_port, Q(31) => NPC_wb_31_port, Q(30) => 
                           NPC_wb_30_port, Q(29) => NPC_wb_29_port, Q(28) => 
                           NPC_wb_28_port, Q(27) => NPC_wb_27_port, Q(26) => 
                           NPC_wb_26_port, Q(25) => NPC_wb_25_port, Q(24) => 
                           NPC_wb_24_port, Q(23) => NPC_wb_23_port, Q(22) => 
                           NPC_wb_22_port, Q(21) => NPC_wb_21_port, Q(20) => 
                           NPC_wb_20_port, Q(19) => NPC_wb_19_port, Q(18) => 
                           NPC_wb_18_port, Q(17) => NPC_wb_17_port, Q(16) => 
                           NPC_wb_16_port, Q(15) => NPC_wb_15_port, Q(14) => 
                           NPC_wb_14_port, Q(13) => NPC_wb_13_port, Q(12) => 
                           NPC_wb_12_port, Q(11) => NPC_wb_11_port, Q(10) => 
                           NPC_wb_10_port, Q(9) => NPC_wb_9_port, Q(8) => 
                           NPC_wb_8_port, Q(7) => NPC_wb_7_port, Q(6) => 
                           NPC_wb_6_port, Q(5) => NPC_wb_5_port, Q(4) => 
                           NPC_wb_4_port, Q(3) => NPC_wb_3_port, Q(2) => 
                           NPC_wb_2_port, Q(1) => NPC_wb_1_port, Q(0) => 
                           NPC_wb_0_port);
   MUX_WB : MUX21_GENERIC_NBIT32_2 port map( A(31) => ALU_wb_31_port, A(30) => 
                           ALU_wb_30_port, A(29) => ALU_wb_29_port, A(28) => 
                           ALU_wb_28_port, A(27) => ALU_wb_27_port, A(26) => 
                           ALU_wb_26_port, A(25) => ALU_wb_25_port, A(24) => 
                           ALU_wb_24_port, A(23) => ALU_wb_23_port, A(22) => 
                           ALU_wb_22_port, A(21) => ALU_wb_21_port, A(20) => 
                           ALU_wb_20_port, A(19) => ALU_wb_19_port, A(18) => 
                           ALU_wb_18_port, A(17) => ALU_wb_17_port, A(16) => 
                           ALU_wb_16_port, A(15) => ALU_wb_15_port, A(14) => 
                           ALU_wb_14_port, A(13) => ALU_wb_13_port, A(12) => 
                           ALU_wb_12_port, A(11) => ALU_wb_11_port, A(10) => 
                           ALU_wb_10_port, A(9) => ALU_wb_9_port, A(8) => 
                           ALU_wb_8_port, A(7) => ALU_wb_7_port, A(6) => 
                           ALU_wb_6_port, A(5) => ALU_wb_5_port, A(4) => 
                           ALU_wb_4_port, A(3) => ALU_wb_3_port, A(2) => 
                           ALU_wb_2_port, A(1) => ALU_wb_1_port, A(0) => 
                           ALU_wb_0_port, B(31) => LMD_wb_31_port, B(30) => 
                           LMD_wb_30_port, B(29) => LMD_wb_29_port, B(28) => 
                           LMD_wb_28_port, B(27) => LMD_wb_27_port, B(26) => 
                           LMD_wb_26_port, B(25) => LMD_wb_25_port, B(24) => 
                           LMD_wb_24_port, B(23) => LMD_wb_23_port, B(22) => 
                           LMD_wb_22_port, B(21) => LMD_wb_21_port, B(20) => 
                           LMD_wb_20_port, B(19) => LMD_wb_19_port, B(18) => 
                           LMD_wb_18_port, B(17) => LMD_wb_17_port, B(16) => 
                           LMD_wb_16_port, B(15) => LMD_wb_15_port, B(14) => 
                           LMD_wb_14_port, B(13) => LMD_wb_13_port, B(12) => 
                           LMD_wb_12_port, B(11) => LMD_wb_11_port, B(10) => 
                           LMD_wb_10_port, B(9) => LMD_wb_9_port, B(8) => 
                           LMD_wb_8_port, B(7) => LMD_wb_7_port, B(6) => 
                           LMD_wb_6_port, B(5) => LMD_wb_5_port, B(4) => 
                           LMD_wb_4_port, B(3) => LMD_wb_3_port, B(2) => 
                           LMD_wb_2_port, B(1) => LMD_wb_1_port, B(0) => 
                           LMD_wb_0_port, SEL => S3, Y(31) => OUT_data_31_port,
                           Y(30) => OUT_data_30_port, Y(29) => OUT_data_29_port
                           , Y(28) => OUT_data_28_port, Y(27) => 
                           OUT_data_27_port, Y(26) => OUT_data_26_port, Y(25) 
                           => OUT_data_25_port, Y(24) => OUT_data_24_port, 
                           Y(23) => OUT_data_23_port, Y(22) => OUT_data_22_port
                           , Y(21) => OUT_data_21_port, Y(20) => 
                           OUT_data_20_port, Y(19) => OUT_data_19_port, Y(18) 
                           => OUT_data_18_port, Y(17) => OUT_data_17_port, 
                           Y(16) => OUT_data_16_port, Y(15) => OUT_data_15_port
                           , Y(14) => OUT_data_14_port, Y(13) => 
                           OUT_data_13_port, Y(12) => OUT_data_12_port, Y(11) 
                           => OUT_data_11_port, Y(10) => OUT_data_10_port, Y(9)
                           => OUT_data_9_port, Y(8) => OUT_data_8_port, Y(7) =>
                           OUT_data_7_port, Y(6) => OUT_data_6_port, Y(5) => 
                           OUT_data_5_port, Y(4) => OUT_data_4_port, Y(3) => 
                           OUT_data_3_port, Y(2) => OUT_data_2_port, Y(1) => 
                           OUT_data_1_port, Y(0) => OUT_data_0_port);
   MUX_jal : MUX21_GENERIC_NBIT32_1 port map( A(31) => NPC_wb_31_port, A(30) =>
                           NPC_wb_30_port, A(29) => NPC_wb_29_port, A(28) => 
                           NPC_wb_28_port, A(27) => NPC_wb_27_port, A(26) => 
                           NPC_wb_26_port, A(25) => NPC_wb_25_port, A(24) => 
                           NPC_wb_24_port, A(23) => NPC_wb_23_port, A(22) => 
                           NPC_wb_22_port, A(21) => NPC_wb_21_port, A(20) => 
                           NPC_wb_20_port, A(19) => NPC_wb_19_port, A(18) => 
                           NPC_wb_18_port, A(17) => NPC_wb_17_port, A(16) => 
                           NPC_wb_16_port, A(15) => NPC_wb_15_port, A(14) => 
                           NPC_wb_14_port, A(13) => NPC_wb_13_port, A(12) => 
                           NPC_wb_12_port, A(11) => NPC_wb_11_port, A(10) => 
                           NPC_wb_10_port, A(9) => NPC_wb_9_port, A(8) => 
                           NPC_wb_8_port, A(7) => NPC_wb_7_port, A(6) => 
                           NPC_wb_6_port, A(5) => NPC_wb_5_port, A(4) => 
                           NPC_wb_4_port, A(3) => NPC_wb_3_port, A(2) => 
                           NPC_wb_2_port, A(1) => NPC_wb_1_port, A(0) => 
                           NPC_wb_0_port, B(31) => OUT_data_31_port, B(30) => 
                           OUT_data_30_port, B(29) => OUT_data_29_port, B(28) 
                           => OUT_data_28_port, B(27) => OUT_data_27_port, 
                           B(26) => OUT_data_26_port, B(25) => OUT_data_25_port
                           , B(24) => OUT_data_24_port, B(23) => 
                           OUT_data_23_port, B(22) => OUT_data_22_port, B(21) 
                           => OUT_data_21_port, B(20) => OUT_data_20_port, 
                           B(19) => OUT_data_19_port, B(18) => OUT_data_18_port
                           , B(17) => OUT_data_17_port, B(16) => 
                           OUT_data_16_port, B(15) => OUT_data_15_port, B(14) 
                           => OUT_data_14_port, B(13) => OUT_data_13_port, 
                           B(12) => OUT_data_12_port, B(11) => OUT_data_11_port
                           , B(10) => OUT_data_10_port, B(9) => OUT_data_9_port
                           , B(8) => OUT_data_8_port, B(7) => OUT_data_7_port, 
                           B(6) => OUT_data_6_port, B(5) => OUT_data_5_port, 
                           B(4) => OUT_data_4_port, B(3) => OUT_data_3_port, 
                           B(2) => OUT_data_2_port, B(1) => OUT_data_1_port, 
                           B(0) => OUT_data_0_port, SEL => sel_saved_reg_wb, 
                           Y(31) => OUT_wb_31_port, Y(30) => OUT_wb_30_port, 
                           Y(29) => OUT_wb_29_port, Y(28) => OUT_wb_28_port, 
                           Y(27) => OUT_wb_27_port, Y(26) => OUT_wb_26_port, 
                           Y(25) => OUT_wb_25_port, Y(24) => OUT_wb_24_port, 
                           Y(23) => OUT_wb_23_port, Y(22) => OUT_wb_22_port, 
                           Y(21) => OUT_wb_21_port, Y(20) => OUT_wb_20_port, 
                           Y(19) => OUT_wb_19_port, Y(18) => OUT_wb_18_port, 
                           Y(17) => OUT_wb_17_port, Y(16) => OUT_wb_16_port, 
                           Y(15) => OUT_wb_15_port, Y(14) => OUT_wb_14_port, 
                           Y(13) => OUT_wb_13_port, Y(12) => OUT_wb_12_port, 
                           Y(11) => OUT_wb_11_port, Y(10) => OUT_wb_10_port, 
                           Y(9) => OUT_wb_9_port, Y(8) => OUT_wb_8_port, Y(7) 
                           => OUT_wb_7_port, Y(6) => OUT_wb_6_port, Y(5) => 
                           OUT_wb_5_port, Y(4) => OUT_wb_4_port, Y(3) => 
                           OUT_wb_3_port, Y(2) => OUT_wb_2_port, Y(1) => 
                           OUT_wb_1_port, Y(0) => OUT_wb_0_port);
   add_256 : DATAPTH_NBIT32_REG_BIT5_DW01_inc_0 port map( A(31) => 
                           PC_fetch0_31_port, A(30) => PC_fetch0_30_port, A(29)
                           => PC_fetch0_29_port, A(28) => PC_fetch0_28_port, 
                           A(27) => PC_fetch0_27_port, A(26) => 
                           PC_fetch0_26_port, A(25) => PC_fetch0_25_port, A(24)
                           => PC_fetch0_24_port, A(23) => PC_fetch0_23_port, 
                           A(22) => PC_fetch0_22_port, A(21) => 
                           PC_fetch0_21_port, A(20) => PC_fetch0_20_port, A(19)
                           => PC_fetch0_19_port, A(18) => PC_fetch0_18_port, 
                           A(17) => PC_fetch0_17_port, A(16) => 
                           PC_fetch0_16_port, A(15) => PC_fetch0_15_port, A(14)
                           => PC_fetch0_14_port, A(13) => PC_fetch0_13_port, 
                           A(12) => PC_fetch0_12_port, A(11) => 
                           PC_fetch0_11_port, A(10) => PC_fetch0_10_port, A(9) 
                           => PC_fetch0_9_port, A(8) => PC_fetch0_8_port, A(7) 
                           => PC_fetch0_7_port, A(6) => PC_fetch0_6_port, A(5) 
                           => PC_fetch0_5_port, A(4) => PC_fetch0_4_port, A(3) 
                           => PC_fetch0_3_port, A(2) => PC_fetch0_2_port, A(1) 
                           => PC_fetch0_1_port, A(0) => PC_fetch0_0_port, 
                           SUM(31) => NPC_31_port, SUM(30) => NPC_30_port, 
                           SUM(29) => NPC_29_port, SUM(28) => NPC_28_port, 
                           SUM(27) => NPC_27_port, SUM(26) => NPC_26_port, 
                           SUM(25) => NPC_25_port, SUM(24) => NPC_24_port, 
                           SUM(23) => NPC_23_port, SUM(22) => NPC_22_port, 
                           SUM(21) => NPC_21_port, SUM(20) => NPC_20_port, 
                           SUM(19) => NPC_19_port, SUM(18) => NPC_18_port, 
                           SUM(17) => NPC_17_port, SUM(16) => NPC_16_port, 
                           SUM(15) => NPC_15_port, SUM(14) => NPC_14_port, 
                           SUM(13) => NPC_13_port, SUM(12) => NPC_12_port, 
                           SUM(11) => NPC_11_port, SUM(10) => NPC_10_port, 
                           SUM(9) => NPC_9_port, SUM(8) => NPC_8_port, SUM(7) 
                           => NPC_7_port, SUM(6) => NPC_6_port, SUM(5) => 
                           NPC_5_port, SUM(4) => NPC_4_port, SUM(3) => 
                           NPC_3_port, SUM(2) => NPC_2_port, SUM(1) => 
                           NPC_1_port, SUM(0) => NPC_0_port);
   U3 : INV_X1 port map( A => n14, ZN => n1);
   U4 : CLKBUF_X1 port map( A => IR_Dec_29_port, Z => n2);
   U5 : BUF_X2 port map( A => RST, Z => n9);
   U6 : BUF_X2 port map( A => RST, Z => n8);
   U7 : BUF_X1 port map( A => n61, Z => n3);
   U8 : BUF_X1 port map( A => n61, Z => n4);
   U9 : BUF_X1 port map( A => N13, Z => n6);
   U10 : BUF_X1 port map( A => N13, Z => n5);
   U11 : BUF_X1 port map( A => N13, Z => n7);
   U12 : NOR4_X1 port map( A1 => IR_Dec_21_port, A2 => IR_Dec_20_port, A3 => 
                           IR_Dec_1_port, A4 => IR_Dec_19_port, ZN => n34);
   U13 : NOR4_X1 port map( A1 => IR_Dec_2_port, A2 => IR_Dec_28_port, A3 => 
                           IR_Dec_26_port, A4 => IR_Dec_25_port, ZN => n36);
   U14 : NAND4_X1 port map( A1 => n35, A2 => n36, A3 => n37, A4 => n38, ZN => 
                           n29);
   U15 : NOR3_X1 port map( A1 => IR_Dec_22_port, A2 => IR_Dec_24_port, A3 => 
                           IR_Dec_23_port, ZN => n35);
   U16 : NOR3_X1 port map( A1 => IR_Dec_3_port, A2 => IR_Dec_5_port, A3 => 
                           IR_Dec_4_port, ZN => n37);
   U17 : NOR4_X1 port map( A1 => IR_Dec_9_port, A2 => IR_Dec_8_port, A3 => 
                           IR_Dec_7_port, A4 => IR_Dec_6_port, ZN => n38);
   U18 : NAND4_X1 port map( A1 => n31, A2 => n32, A3 => n33, A4 => n34, ZN => 
                           n30);
   U19 : NOR3_X1 port map( A1 => IR_Dec_0_port, A2 => IR_Dec_11_port, A3 => 
                           IR_Dec_10_port, ZN => n31);
   U20 : NOR3_X1 port map( A1 => IR_Dec_16_port, A2 => IR_Dec_18_port, A3 => 
                           IR_Dec_17_port, ZN => n33);
   U21 : NOR4_X1 port map( A1 => IR_Dec_15_port, A2 => IR_Dec_14_port, A3 => 
                           IR_Dec_13_port, A4 => IR_Dec_12_port, ZN => n32);
   U22 : INV_X1 port map( A => n23, ZN => n12);
   U23 : INV_X1 port map( A => IR_Dec_31_port, ZN => n13_port);
   U24 : INV_X1 port map( A => IR_Dec_28_port, ZN => n16);
   U25 : INV_X1 port map( A => n26, ZN => n15);
   U26 : AOI21_X1 port map( B1 => n27, B2 => n28, A => IR_Dec_27_port, ZN => 
                           n26);
   U27 : OAI21_X1 port map( B1 => n16, B2 => IR_Dec_26_port, A => n1, ZN => n28
                           );
   U28 : OR2_X1 port map( A1 => n29, A2 => n30, ZN => n27);
   U29 : AOI21_X1 port map( B1 => jump_en, B2 => n21, A => n11, ZN => 
                           wr_signal_mem1);
   U30 : NAND4_X1 port map( A1 => IR_26_mem_1_port, A2 => IR_26_mem_0_port, A3 
                           => n22, A4 => n10, ZN => n21);
   U31 : INV_X1 port map( A => wr_signal_mem, ZN => n11);
   U32 : INV_X1 port map( A => IR_26_mem_2_port, ZN => n10);
   U33 : INV_X1 port map( A => IR_Dec_30_port, ZN => n14);
   U34 : NAND4_X1 port map( A1 => IR_26_mem_2_port, A2 => IR_26_mem_0_port, A3 
                           => IR_26_mem_4_port, A4 => n39, ZN => N13);
   U35 : NOR3_X1 port map( A1 => IR_26_mem_1_port, A2 => IR_26_mem_5_port, A3 
                           => IR_26_mem_3_port, ZN => n39);
   U36 : AOI22_X1 port map( A1 => n51, A2 => instruction_alu(4), B1 => 
                           instruction_alu(3), B2 => n59, ZN => n50);
   U37 : INV_X1 port map( A => instruction_alu(4), ZN => n59);
   U38 : NOR2_X1 port map( A1 => instruction_alu(3), A2 => n60, ZN => n51);
   U39 : OR2_X1 port map( A1 => cond_mem, A2 => jump_en, ZN => sel_npc);
   U40 : INV_X1 port map( A => instruction_alu(5), ZN => n60);
   U41 : INV_X1 port map( A => sb_op, ZN => n61);
   U42 : INV_X1 port map( A => instruction_alu(2), ZN => n58);
   U43 : NOR2_X1 port map( A1 => IR_26_mem_5_port, A2 => IR_26_mem_3_port, ZN 
                           => n22);
   U44 : OR4_X1 port map( A1 => n48, A2 => n49, A3 => WM, A4 => RM, ZN => 
                           DATA_MEM_ENABLE);
   U45 : NOR4_X1 port map( A1 => instruction_alu(1), A2 => n50, A3 => n58, A4 
                           => n57, ZN => n49);
   U46 : NOR4_X1 port map( A1 => n52, A2 => n60, A3 => instruction_alu(0), A4 
                           => instruction_alu(2), ZN => n48);
   U47 : INV_X1 port map( A => instruction_alu(0), ZN => n57);
   U48 : AND2_X1 port map( A1 => IR_26_mem_0_port, A2 => jump_en, ZN => 
                           sel_saved_reg);
   U49 : INV_X1 port map( A => n41, ZN => DATA_MEM_IN(6));
   U50 : AOI22_X1 port map( A1 => n3, A2 => regB_mem_6_port, B1 => sb_op, B2 =>
                           regB_mem_30_port, ZN => n41);
   U51 : INV_X1 port map( A => n42, ZN => DATA_MEM_IN(5));
   U52 : AOI22_X1 port map( A1 => n3, A2 => regB_mem_5_port, B1 => sb_op, B2 =>
                           regB_mem_29_port, ZN => n42);
   U53 : INV_X1 port map( A => n43, ZN => DATA_MEM_IN(4));
   U54 : AOI22_X1 port map( A1 => n3, A2 => regB_mem_4_port, B1 => sb_op, B2 =>
                           regB_mem_28_port, ZN => n43);
   U55 : INV_X1 port map( A => n44, ZN => DATA_MEM_IN(3));
   U56 : AOI22_X1 port map( A1 => n3, A2 => regB_mem_3_port, B1 => sb_op, B2 =>
                           regB_mem_27_port, ZN => n44);
   U57 : INV_X1 port map( A => n45, ZN => DATA_MEM_IN(2));
   U58 : AOI22_X1 port map( A1 => n3, A2 => regB_mem_2_port, B1 => sb_op, B2 =>
                           regB_mem_26_port, ZN => n45);
   U59 : INV_X1 port map( A => n46, ZN => DATA_MEM_IN(1));
   U60 : AOI22_X1 port map( A1 => sb_op, A2 => regB_mem_25_port, B1 => n3, B2 
                           => regB_mem_1_port, ZN => n46);
   U61 : INV_X1 port map( A => n47, ZN => DATA_MEM_IN(0));
   U62 : AOI22_X1 port map( A1 => sb_op, A2 => regB_mem_24_port, B1 => n3, B2 
                           => regB_mem_0_port, ZN => n47);
   U63 : INV_X1 port map( A => n40, ZN => DATA_MEM_IN(7));
   U64 : AOI22_X1 port map( A1 => n3, A2 => regB_mem_7_port, B1 => 
                           regB_mem_31_port, B2 => sb_op, ZN => n40);
   U65 : AND2_X1 port map( A1 => n4, A2 => regB_mem_31_port, ZN => 
                           DATA_MEM_IN(31));
   U66 : AND2_X1 port map( A1 => n4, A2 => regB_mem_30_port, ZN => 
                           DATA_MEM_IN(30));
   U67 : AND2_X1 port map( A1 => n4, A2 => regB_mem_29_port, ZN => 
                           DATA_MEM_IN(29));
   U68 : AND2_X1 port map( A1 => n4, A2 => regB_mem_28_port, ZN => 
                           DATA_MEM_IN(28));
   U69 : AND2_X1 port map( A1 => n4, A2 => regB_mem_27_port, ZN => 
                           DATA_MEM_IN(27));
   U70 : AND2_X1 port map( A1 => n4, A2 => regB_mem_26_port, ZN => 
                           DATA_MEM_IN(26));
   U71 : AND2_X1 port map( A1 => n4, A2 => regB_mem_25_port, ZN => 
                           DATA_MEM_IN(25));
   U72 : AND2_X1 port map( A1 => n4, A2 => regB_mem_24_port, ZN => 
                           DATA_MEM_IN(24));
   U73 : AND2_X1 port map( A1 => regB_mem_14_port, A2 => n3, ZN => 
                           DATA_MEM_IN(14));
   U74 : AND2_X1 port map( A1 => regB_mem_13_port, A2 => n3, ZN => 
                           DATA_MEM_IN(13));
   U75 : AND2_X1 port map( A1 => regB_mem_12_port, A2 => n3, ZN => 
                           DATA_MEM_IN(12));
   U76 : AND2_X1 port map( A1 => regB_mem_11_port, A2 => n3, ZN => 
                           DATA_MEM_IN(11));
   U77 : AND2_X1 port map( A1 => regB_mem_10_port, A2 => n3, ZN => 
                           DATA_MEM_IN(10));
   U78 : AND2_X1 port map( A1 => regB_mem_9_port, A2 => n3, ZN => 
                           DATA_MEM_IN(9));
   U79 : AND2_X1 port map( A1 => regB_mem_23_port, A2 => n4, ZN => 
                           DATA_MEM_IN(23));
   U84 : AND2_X1 port map( A1 => regB_mem_22_port, A2 => n4, ZN => 
                           DATA_MEM_IN(22));
   U85 : AND2_X1 port map( A1 => regB_mem_21_port, A2 => n4, ZN => 
                           DATA_MEM_IN(21));
   U86 : AND2_X1 port map( A1 => regB_mem_20_port, A2 => n4, ZN => 
                           DATA_MEM_IN(20));
   U87 : AND2_X1 port map( A1 => regB_mem_19_port, A2 => n4, ZN => 
                           DATA_MEM_IN(19));
   U88 : AND2_X1 port map( A1 => regB_mem_18_port, A2 => n4, ZN => 
                           DATA_MEM_IN(18));
   U89 : AND2_X1 port map( A1 => regB_mem_17_port, A2 => n4, ZN => 
                           DATA_MEM_IN(17));
   U90 : AND2_X1 port map( A1 => regB_mem_16_port, A2 => n4, ZN => 
                           DATA_MEM_IN(16));
   U91 : AND2_X1 port map( A1 => regB_mem_15_port, A2 => n4, ZN => 
                           DATA_MEM_IN(15));
   U92 : AND2_X1 port map( A1 => regB_mem_8_port, A2 => n4, ZN => 
                           DATA_MEM_IN(8));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity 
   dlx_cu_MICROCODE_MEM_SIZE62_FUNC_SIZE11_OP_CODE_SIZE6_IR_SIZE32_CW_SIZE15 is

   port( Clk, Rst : in std_logic;  IR_IN : in std_logic_vector (31 downto 0);  
         IR_LATCH_EN, NPC_LATCH_EN, RegA_LATCH_EN, RegB_LATCH_EN, 
         RegIMM_LATCH_EN, MUXA_SEL, MUXB_SEL, ALU_OUTREG_EN, EQ_COND : out 
         std_logic;  ALU_OPCODE : out std_logic_vector (0 to 5);  
         signed_unsigned, DRAM_WE, LMD_LATCH_EN, JUMP_EN, PC_LATCH_EN, 
         WB_MUX_SEL, RF_WE, lhi_sel, sb_op, s_trap, s_ret : out std_logic);

end dlx_cu_MICROCODE_MEM_SIZE62_FUNC_SIZE11_OP_CODE_SIZE6_IR_SIZE32_CW_SIZE15;

architecture SYN_dlx_cu_hw of 
   dlx_cu_MICROCODE_MEM_SIZE62_FUNC_SIZE11_OP_CODE_SIZE6_IR_SIZE32_CW_SIZE15 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component AND2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X2
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component 
      dlx_cu_MICROCODE_MEM_SIZE62_FUNC_SIZE11_OP_CODE_SIZE6_IR_SIZE32_CW_SIZE15_DW01_inc_5
      port( A : in std_logic_vector (31 downto 0);  SUM : out std_logic_vector 
            (31 downto 0));
   end component;
   
   component 
      dlx_cu_MICROCODE_MEM_SIZE62_FUNC_SIZE11_OP_CODE_SIZE6_IR_SIZE32_CW_SIZE15_DW01_inc_4
      port( A : in std_logic_vector (31 downto 0);  SUM : out std_logic_vector 
            (31 downto 0));
   end component;
   
   component 
      dlx_cu_MICROCODE_MEM_SIZE62_FUNC_SIZE11_OP_CODE_SIZE6_IR_SIZE32_CW_SIZE15_DW01_inc_3
      port( A : in std_logic_vector (31 downto 0);  SUM : out std_logic_vector 
            (31 downto 0));
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal signed_unsigned_port, sb_op_port, aluOpcode1_5_port, 
      aluOpcode1_4_port, aluOpcode1_3_port, aluOpcode1_2_port, 
      aluOpcode1_1_port, aluOpcode1_0_port, aluOpcode2_5_port, 
      aluOpcode2_4_port, aluOpcode2_3_port, aluOpcode2_2_port, 
      aluOpcode2_1_port, aluOpcode2_0_port, iterator_trap_31_port, 
      iterator_trap_30_port, iterator_trap_29_port, iterator_trap_28_port, 
      iterator_trap_27_port, iterator_trap_26_port, iterator_trap_25_port, 
      iterator_trap_24_port, iterator_trap_23_port, iterator_trap_22_port, 
      iterator_trap_21_port, iterator_trap_20_port, iterator_trap_19_port, 
      iterator_trap_18_port, iterator_trap_17_port, iterator_trap_16_port, 
      iterator_trap_15_port, iterator_trap_14_port, iterator_trap_13_port, 
      iterator_trap_12_port, iterator_trap_11_port, iterator_trap_10_port, 
      iterator_trap_9_port, iterator_trap_8_port, iterator_trap_7_port, 
      iterator_trap_6_port, iterator_trap_5_port, iterator_trap_4_port, 
      iterator_trap_3_port, iterator_trap_2_port, iterator_trap_1_port, 
      iterator_trap_0_port, N34, N35, N36, N37, N38, N39, N40, N41, N42, N43, 
      N44, N45, N46, N47, N48, N49, N50, N51, N52, N53, N54, N55, N56, N57, N58
      , N59, N60, N61, N62, N63, N64, N65, iterator_ret_31_port, 
      iterator_ret_30_port, iterator_ret_29_port, iterator_ret_28_port, 
      iterator_ret_27_port, iterator_ret_26_port, iterator_ret_25_port, 
      iterator_ret_24_port, iterator_ret_23_port, iterator_ret_22_port, 
      iterator_ret_21_port, iterator_ret_20_port, iterator_ret_19_port, 
      iterator_ret_18_port, iterator_ret_17_port, iterator_ret_16_port, 
      iterator_ret_15_port, iterator_ret_14_port, iterator_ret_13_port, 
      iterator_ret_12_port, iterator_ret_11_port, iterator_ret_10_port, 
      iterator_ret_9_port, iterator_ret_8_port, iterator_ret_7_port, 
      iterator_ret_6_port, iterator_ret_5_port, iterator_ret_4_port, 
      iterator_ret_3_port, iterator_ret_2_port, iterator_ret_1_port, 
      iterator_ret_0_port, N145, N146, N147, N148, N149, N150, N151, N152, N153
      , N154, N155, N156, N157, N158, N159, N160, N161, N162, N163, N164, N165,
      N166, N167, N168, N169, N170, N171, N172, N173, N174, N175, N176, 
      iterator1_31_port, iterator1_30_port, iterator1_29_port, 
      iterator1_28_port, iterator1_27_port, iterator1_26_port, 
      iterator1_25_port, iterator1_24_port, iterator1_23_port, 
      iterator1_22_port, iterator1_21_port, iterator1_20_port, 
      iterator1_19_port, iterator1_18_port, iterator1_17_port, 
      iterator1_16_port, iterator1_15_port, iterator1_14_port, 
      iterator1_13_port, iterator1_12_port, iterator1_11_port, 
      iterator1_10_port, iterator1_9_port, iterator1_8_port, iterator1_7_port, 
      iterator1_6_port, iterator1_5_port, iterator1_4_port, iterator1_3_port, 
      iterator1_2_port, iterator1_1_port, iterator1_0_port, N253, N254, N255, 
      N256, N257, N258, N259, N260, N261, N262, N263, N264, N265, N266, N267, 
      N268, N269, N270, N271, N272, N273, N274, N275, N276, N277, N278, N279, 
      N280, N281, N282, N283, N284, aluOpcode_i_5_port, aluOpcode_i_4_port, 
      aluOpcode_i_3_port, aluOpcode_i_2_port, aluOpcode_i_1_port, 
      aluOpcode_i_0_port, signed_unsigned_i, N550, N551, n271_port, n272_port, 
      n273_port, n274_port, n275_port, n276_port, n277_port, n278_port, 
      n279_port, n280_port, n281_port, n282_port, n283_port, n284_port, n285, 
      n286, n287, n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, 
      n298, n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309, 
      n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320, n321, 
      n322, n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, 
      n334, n336, n339, n340, n343, n344, n345, n377, n379, n380, n381, n382, 
      n383, n384, n385, n386, n387, n388, n389, n390, n391, n392, n393, n394, 
      n395, n396, n397, n398, n399, n400, n401, n402, n403, n404, n405, n406, 
      n407, n408, n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, 
      n419, n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, 
      n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, 
      n443, n444, n445, n446, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12
      , n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, 
      n27, n28, n29, n30, n31, n32, n33, n34_port, n35_port, n36_port, n37_port
      , n38_port, n39_port, n40_port, n41_port, n42_port, n43_port, n44_port, 
      n45_port, n46_port, n47_port, n48_port, n49_port, n50_port, n51_port, 
      n52_port, n53_port, n54_port, n55_port, n56_port, n57_port, n58_port, 
      n59_port, n60_port, n61_port, n62_port, n63_port, n64_port, n65_port, n66
      , n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, 
      n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95
      , n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, 
      n108, n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119, 
      n120, n121, n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, 
      n132, n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, 
      n144, n145_port, n146_port, n147_port, n148_port, n149_port, n150_port, 
      n151_port, n152_port, n153_port, n154_port, n155_port, n156_port, 
      n157_port, n158_port, n159_port, n160_port, n161_port, n162_port, 
      n163_port, n164_port, n165_port, n166_port, n167_port, n168_port, 
      n169_port, n170_port, n171_port, n172_port, n173_port, n174_port, 
      n175_port, n176_port, n177, n178, n179, n180, n181, n182, n183, n184, 
      n185, n186, n187, n188, n189, n190, n191, n192, n193, n194, n195, n196, 
      n197, n198, n199, n200, n201, n202, n203, n204, n205, n206, n207, n208, 
      n209, n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, 
      n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232, 
      n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243, n244, 
      n245, n246, n247, n248, n249, n250, n251, n252, n253_port, n254_port, 
      n255_port, n256_port, n257_port, n258_port, n259_port, n260_port, 
      n261_port, n262_port, n263_port, n264_port, n265_port, n266_port, 
      n267_port, n268_port, n269_port, n270_port, n335, n337, n338, n341, n342,
      n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, 
      n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369, 
      n370, n371, n372, n373, n374, n375, n376, n378, n447, n448, n449, n450, 
      n451, n452, n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, 
      n463, n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, 
      n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, 
      n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, 
      n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, 
      n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, 
      n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, 
      n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, 
      n547, n548, n549, n_2358, n_2359, n_2360, n_2361, n_2362, n_2363, n_2364,
      n_2365, n_2366, n_2367, n_2368, n_2369, n_2370, n_2371, n_2372, n_2373, 
      n_2374, n_2375, n_2376, n_2377, n_2378, n_2379 : std_logic;

begin
   signed_unsigned <= signed_unsigned_port;
   sb_op <= sb_op_port;
   
   aluOpcode1_reg_5_inst : DFFR_X1 port map( D => aluOpcode_i_5_port, CK => Clk
                           , RN => n64_port, Q => aluOpcode1_5_port, QN => 
                           n_2358);
   aluOpcode1_reg_4_inst : DFFR_X1 port map( D => aluOpcode_i_4_port, CK => Clk
                           , RN => n63_port, Q => aluOpcode1_4_port, QN => 
                           n_2359);
   aluOpcode1_reg_3_inst : DFFR_X1 port map( D => aluOpcode_i_3_port, CK => Clk
                           , RN => n63_port, Q => aluOpcode1_3_port, QN => 
                           n_2360);
   aluOpcode1_reg_2_inst : DFFR_X1 port map( D => aluOpcode_i_2_port, CK => Clk
                           , RN => n63_port, Q => aluOpcode1_2_port, QN => 
                           n_2361);
   aluOpcode1_reg_1_inst : DFFR_X1 port map( D => aluOpcode_i_1_port, CK => Clk
                           , RN => n63_port, Q => aluOpcode1_1_port, QN => 
                           n_2362);
   aluOpcode1_reg_0_inst : DFFR_X1 port map( D => aluOpcode_i_0_port, CK => Clk
                           , RN => n63_port, Q => aluOpcode1_0_port, QN => 
                           n_2363);
   aluOpcode2_reg_5_inst : DFFR_X1 port map( D => aluOpcode1_5_port, CK => Clk,
                           RN => n63_port, Q => aluOpcode2_5_port, QN => n_2364
                           );
   aluOpcode2_reg_4_inst : DFFR_X1 port map( D => aluOpcode1_4_port, CK => Clk,
                           RN => n63_port, Q => aluOpcode2_4_port, QN => n_2365
                           );
   aluOpcode2_reg_3_inst : DFFR_X1 port map( D => aluOpcode1_3_port, CK => Clk,
                           RN => n63_port, Q => aluOpcode2_3_port, QN => n_2366
                           );
   aluOpcode2_reg_2_inst : DFFR_X1 port map( D => aluOpcode1_2_port, CK => Clk,
                           RN => n63_port, Q => aluOpcode2_2_port, QN => n_2367
                           );
   aluOpcode2_reg_1_inst : DFFR_X1 port map( D => aluOpcode1_1_port, CK => Clk,
                           RN => n64_port, Q => aluOpcode2_1_port, QN => n_2368
                           );
   aluOpcode2_reg_0_inst : DFFR_X1 port map( D => aluOpcode1_0_port, CK => Clk,
                           RN => n64_port, Q => aluOpcode2_0_port, QN => n_2369
                           );
   aluOpcode3_reg_5_inst : DFFR_X1 port map( D => aluOpcode2_5_port, CK => Clk,
                           RN => n64_port, Q => ALU_OPCODE(0), QN => n_2370);
   aluOpcode3_reg_4_inst : DFFR_X1 port map( D => aluOpcode2_4_port, CK => Clk,
                           RN => n64_port, Q => ALU_OPCODE(1), QN => n_2371);
   aluOpcode3_reg_3_inst : DFFR_X1 port map( D => aluOpcode2_3_port, CK => Clk,
                           RN => n64_port, Q => ALU_OPCODE(2), QN => n_2372);
   aluOpcode3_reg_2_inst : DFFR_X1 port map( D => aluOpcode2_2_port, CK => Clk,
                           RN => n64_port, Q => ALU_OPCODE(3), QN => n_2373);
   aluOpcode3_reg_1_inst : DFFR_X1 port map( D => aluOpcode2_1_port, CK => Clk,
                           RN => n64_port, Q => ALU_OPCODE(4), QN => n_2374);
   aluOpcode3_reg_0_inst : DFFR_X1 port map( D => aluOpcode2_0_port, CK => Clk,
                           RN => n64_port, Q => ALU_OPCODE(5), QN => n_2375);
   iterator_ret_reg_26_inst : DFF_X1 port map( D => n439, CK => Clk, Q => 
                           iterator_ret_26_port, QN => n329);
   iterator_ret_reg_20_inst : DFF_X1 port map( D => n433, CK => Clk, Q => 
                           iterator_ret_20_port, QN => n323);
   iterator_ret_reg_19_inst : DFF_X1 port map( D => n432, CK => Clk, Q => 
                           iterator_ret_19_port, QN => n322);
   iterator_ret_reg_16_inst : DFF_X1 port map( D => n429, CK => Clk, Q => 
                           iterator_ret_16_port, QN => n319);
   iterator_ret_reg_14_inst : DFF_X1 port map( D => n427, CK => Clk, Q => 
                           iterator_ret_14_port, QN => n317);
   iterator_ret_reg_8_inst : DFF_X1 port map( D => n421, CK => Clk, Q => 
                           iterator_ret_8_port, QN => n311);
   iterator_ret_reg_7_inst : DFF_X1 port map( D => n420, CK => Clk, Q => 
                           iterator_ret_7_port, QN => n310);
   iterator1_reg_30_inst : DFF_X1 port map( D => n519, CK => Clk, Q => 
                           iterator1_30_port, QN => n133);
   iterator1_reg_29_inst : DFF_X1 port map( D => n520, CK => Clk, Q => 
                           iterator1_29_port, QN => n131);
   iterator1_reg_28_inst : DFF_X1 port map( D => n521, CK => Clk, Q => 
                           iterator1_28_port, QN => n129);
   iterator1_reg_27_inst : DFF_X1 port map( D => n522, CK => Clk, Q => 
                           iterator1_27_port, QN => n127);
   iterator1_reg_26_inst : DFF_X1 port map( D => n523, CK => Clk, Q => 
                           iterator1_26_port, QN => n125);
   iterator1_reg_25_inst : DFF_X1 port map( D => n524, CK => Clk, Q => 
                           iterator1_25_port, QN => n123);
   iterator1_reg_24_inst : DFF_X1 port map( D => n525, CK => Clk, Q => 
                           iterator1_24_port, QN => n121);
   iterator1_reg_23_inst : DFF_X1 port map( D => n526, CK => Clk, Q => 
                           iterator1_23_port, QN => n119);
   iterator1_reg_22_inst : DFF_X1 port map( D => n527, CK => Clk, Q => 
                           iterator1_22_port, QN => n117);
   iterator1_reg_21_inst : DFF_X1 port map( D => n528, CK => Clk, Q => 
                           iterator1_21_port, QN => n115);
   iterator1_reg_20_inst : DFF_X1 port map( D => n529, CK => Clk, Q => 
                           iterator1_20_port, QN => n113);
   iterator1_reg_19_inst : DFF_X1 port map( D => n530, CK => Clk, Q => 
                           iterator1_19_port, QN => n111);
   iterator1_reg_18_inst : DFF_X1 port map( D => n531, CK => Clk, Q => 
                           iterator1_18_port, QN => n109);
   iterator1_reg_17_inst : DFF_X1 port map( D => n532, CK => Clk, Q => 
                           iterator1_17_port, QN => n107);
   iterator1_reg_16_inst : DFF_X1 port map( D => n533, CK => Clk, Q => 
                           iterator1_16_port, QN => n105);
   iterator1_reg_15_inst : DFF_X1 port map( D => n534, CK => Clk, Q => 
                           iterator1_15_port, QN => n103);
   iterator1_reg_14_inst : DFF_X1 port map( D => n535, CK => Clk, Q => 
                           iterator1_14_port, QN => n101);
   iterator1_reg_13_inst : DFF_X1 port map( D => n536, CK => Clk, Q => 
                           iterator1_13_port, QN => n99);
   iterator1_reg_12_inst : DFF_X1 port map( D => n537, CK => Clk, Q => 
                           iterator1_12_port, QN => n97);
   iterator1_reg_11_inst : DFF_X1 port map( D => n538, CK => Clk, Q => 
                           iterator1_11_port, QN => n95);
   iterator1_reg_10_inst : DFF_X1 port map( D => n539, CK => Clk, Q => 
                           iterator1_10_port, QN => n93);
   iterator1_reg_9_inst : DFF_X1 port map( D => n540, CK => Clk, Q => 
                           iterator1_9_port, QN => n91);
   iterator1_reg_8_inst : DFF_X1 port map( D => n541, CK => Clk, Q => 
                           iterator1_8_port, QN => n89);
   iterator1_reg_7_inst : DFF_X1 port map( D => n542, CK => Clk, Q => 
                           iterator1_7_port, QN => n87);
   iterator1_reg_6_inst : DFF_X1 port map( D => n543, CK => Clk, Q => 
                           iterator1_6_port, QN => n85);
   iterator1_reg_5_inst : DFF_X1 port map( D => n544, CK => Clk, Q => 
                           iterator1_5_port, QN => n83);
   iterator1_reg_4_inst : DFF_X1 port map( D => n545, CK => Clk, Q => 
                           iterator1_4_port, QN => n81);
   iterator1_reg_31_inst : DFF_X1 port map( D => n549, CK => Clk, Q => 
                           iterator1_31_port, QN => n76);
   sb_op_reg : DFF_X1 port map( D => n345, CK => Clk, Q => sb_op_port, QN => 
                           n_2376);
   signed_unsigned_i_reg : DLH_X1 port map( G => N550, D => N551, Q => 
                           signed_unsigned_i);
   signed_unsigned_1_reg : DFF_X1 port map( D => n344, CK => Clk, Q => n249, QN
                           => n_2377);
   signed_unsigned_2_reg : DFF_X1 port map( D => n343, CK => Clk, Q => 
                           signed_unsigned_port, QN => n_2378);
   RF_WE <= '0';
   WB_MUX_SEL <= '0';
   PC_LATCH_EN <= '0';
   JUMP_EN <= '0';
   LMD_LATCH_EN <= '0';
   DRAM_WE <= '0';
   EQ_COND <= '0';
   ALU_OUTREG_EN <= '0';
   MUXB_SEL <= '0';
   MUXA_SEL <= '0';
   RegIMM_LATCH_EN <= '0';
   RegB_LATCH_EN <= '0';
   RegA_LATCH_EN <= '0';
   NPC_LATCH_EN <= '0';
   IR_LATCH_EN <= '0';
   add_239 : 
                           dlx_cu_MICROCODE_MEM_SIZE62_FUNC_SIZE11_OP_CODE_SIZE6_IR_SIZE32_CW_SIZE15_DW01_inc_3 
                           port map( A(31) => iterator_ret_31_port, A(30) => 
                           iterator_ret_30_port, A(29) => iterator_ret_29_port,
                           A(28) => iterator_ret_28_port, A(27) => 
                           iterator_ret_27_port, A(26) => iterator_ret_26_port,
                           A(25) => iterator_ret_25_port, A(24) => 
                           iterator_ret_24_port, A(23) => iterator_ret_23_port,
                           A(22) => iterator_ret_22_port, A(21) => 
                           iterator_ret_21_port, A(20) => iterator_ret_20_port,
                           A(19) => iterator_ret_19_port, A(18) => 
                           iterator_ret_18_port, A(17) => iterator_ret_17_port,
                           A(16) => iterator_ret_16_port, A(15) => 
                           iterator_ret_15_port, A(14) => iterator_ret_14_port,
                           A(13) => iterator_ret_13_port, A(12) => 
                           iterator_ret_12_port, A(11) => iterator_ret_11_port,
                           A(10) => iterator_ret_10_port, A(9) => 
                           iterator_ret_9_port, A(8) => iterator_ret_8_port, 
                           A(7) => iterator_ret_7_port, A(6) => 
                           iterator_ret_6_port, A(5) => iterator_ret_5_port, 
                           A(4) => iterator_ret_4_port, A(3) => 
                           iterator_ret_3_port, A(2) => iterator_ret_2_port, 
                           A(1) => iterator_ret_1_port, A(0) => 
                           iterator_ret_0_port, SUM(31) => N176, SUM(30) => 
                           N175, SUM(29) => N174, SUM(28) => N173, SUM(27) => 
                           N172, SUM(26) => N171, SUM(25) => N170, SUM(24) => 
                           N169, SUM(23) => N168, SUM(22) => N167, SUM(21) => 
                           N166, SUM(20) => N165, SUM(19) => N164, SUM(18) => 
                           N163, SUM(17) => N162, SUM(16) => N161, SUM(15) => 
                           N160, SUM(14) => N159, SUM(13) => N158, SUM(12) => 
                           N157, SUM(11) => N156, SUM(10) => N155, SUM(9) => 
                           N154, SUM(8) => N153, SUM(7) => N152, SUM(6) => N151
                           , SUM(5) => N150, SUM(4) => N149, SUM(3) => N148, 
                           SUM(2) => N147, SUM(1) => N146, SUM(0) => N145);
   add_217 : 
                           dlx_cu_MICROCODE_MEM_SIZE62_FUNC_SIZE11_OP_CODE_SIZE6_IR_SIZE32_CW_SIZE15_DW01_inc_4 
                           port map( A(31) => iterator_trap_31_port, A(30) => 
                           iterator_trap_30_port, A(29) => 
                           iterator_trap_29_port, A(28) => 
                           iterator_trap_28_port, A(27) => 
                           iterator_trap_27_port, A(26) => 
                           iterator_trap_26_port, A(25) => 
                           iterator_trap_25_port, A(24) => 
                           iterator_trap_24_port, A(23) => 
                           iterator_trap_23_port, A(22) => 
                           iterator_trap_22_port, A(21) => 
                           iterator_trap_21_port, A(20) => 
                           iterator_trap_20_port, A(19) => 
                           iterator_trap_19_port, A(18) => 
                           iterator_trap_18_port, A(17) => 
                           iterator_trap_17_port, A(16) => 
                           iterator_trap_16_port, A(15) => 
                           iterator_trap_15_port, A(14) => 
                           iterator_trap_14_port, A(13) => 
                           iterator_trap_13_port, A(12) => 
                           iterator_trap_12_port, A(11) => 
                           iterator_trap_11_port, A(10) => 
                           iterator_trap_10_port, A(9) => iterator_trap_9_port,
                           A(8) => iterator_trap_8_port, A(7) => 
                           iterator_trap_7_port, A(6) => iterator_trap_6_port, 
                           A(5) => iterator_trap_5_port, A(4) => 
                           iterator_trap_4_port, A(3) => iterator_trap_3_port, 
                           A(2) => iterator_trap_2_port, A(1) => 
                           iterator_trap_1_port, A(0) => iterator_trap_0_port, 
                           SUM(31) => N65, SUM(30) => N64, SUM(29) => N63, 
                           SUM(28) => N62, SUM(27) => N61, SUM(26) => N60, 
                           SUM(25) => N59, SUM(24) => N58, SUM(23) => N57, 
                           SUM(22) => N56, SUM(21) => N55, SUM(20) => N54, 
                           SUM(19) => N53, SUM(18) => N52, SUM(17) => N51, 
                           SUM(16) => N50, SUM(15) => N49, SUM(14) => N48, 
                           SUM(13) => N47, SUM(12) => N46, SUM(11) => N45, 
                           SUM(10) => N44, SUM(9) => N43, SUM(8) => N42, SUM(7)
                           => N41, SUM(6) => N40, SUM(5) => N39, SUM(4) => N38,
                           SUM(3) => N37, SUM(2) => N36, SUM(1) => N35, SUM(0) 
                           => N34);
   add_258 : 
                           dlx_cu_MICROCODE_MEM_SIZE62_FUNC_SIZE11_OP_CODE_SIZE6_IR_SIZE32_CW_SIZE15_DW01_inc_5 
                           port map( A(31) => iterator1_31_port, A(30) => 
                           iterator1_30_port, A(29) => iterator1_29_port, A(28)
                           => iterator1_28_port, A(27) => iterator1_27_port, 
                           A(26) => iterator1_26_port, A(25) => 
                           iterator1_25_port, A(24) => iterator1_24_port, A(23)
                           => iterator1_23_port, A(22) => iterator1_22_port, 
                           A(21) => iterator1_21_port, A(20) => 
                           iterator1_20_port, A(19) => iterator1_19_port, A(18)
                           => iterator1_18_port, A(17) => iterator1_17_port, 
                           A(16) => iterator1_16_port, A(15) => 
                           iterator1_15_port, A(14) => iterator1_14_port, A(13)
                           => iterator1_13_port, A(12) => iterator1_12_port, 
                           A(11) => iterator1_11_port, A(10) => 
                           iterator1_10_port, A(9) => iterator1_9_port, A(8) =>
                           iterator1_8_port, A(7) => iterator1_7_port, A(6) => 
                           iterator1_6_port, A(5) => iterator1_5_port, A(4) => 
                           iterator1_4_port, A(3) => iterator1_3_port, A(2) => 
                           iterator1_2_port, A(1) => iterator1_1_port, A(0) => 
                           iterator1_0_port, SUM(31) => N284, SUM(30) => N283, 
                           SUM(29) => N282, SUM(28) => N281, SUM(27) => N280, 
                           SUM(26) => N279, SUM(25) => N278, SUM(24) => N277, 
                           SUM(23) => N276, SUM(22) => N275, SUM(21) => N274, 
                           SUM(20) => N273, SUM(19) => N272, SUM(18) => N271, 
                           SUM(17) => N270, SUM(16) => N269, SUM(15) => N268, 
                           SUM(14) => N267, SUM(13) => N266, SUM(12) => N265, 
                           SUM(11) => N264, SUM(10) => N263, SUM(9) => N262, 
                           SUM(8) => N261, SUM(7) => N260, SUM(6) => N259, 
                           SUM(5) => N258, SUM(4) => N257, SUM(3) => N256, 
                           SUM(2) => N255, SUM(1) => N254, SUM(0) => N253);
   iterator_ret_reg_21_inst : DFF_X1 port map( D => n434, CK => Clk, Q => 
                           iterator_ret_21_port, QN => n324);
   iterator_ret_reg_24_inst : DFF_X1 port map( D => n437, CK => Clk, Q => 
                           iterator_ret_24_port, QN => n327);
   lhi_sel_reg : DFF_X1 port map( D => n377, CK => Clk, Q => lhi_sel, QN => 
                           n336);
   iterator1_reg_3_inst : DFF_X1 port map( D => n546, CK => Clk, Q => 
                           iterator1_3_port, QN => n40_port);
   iterator1_reg_2_inst : DFF_X1 port map( D => n547, CK => Clk, Q => 
                           iterator1_2_port, QN => n41_port);
   iterator1_reg_1_inst : DFF_X1 port map( D => n548, CK => Clk, Q => 
                           iterator1_1_port, QN => n42_port);
   iterator1_reg_0_inst : DFF_X1 port map( D => n518, CK => Clk, Q => 
                           iterator1_0_port, QN => n43_port);
   s_ret_reg : DFF_X1 port map( D => n379, CK => Clk, Q => s_ret, QN => n340);
   iterator_trap_reg_0_inst : DFF_X1 port map( D => n381, CK => Clk, Q => 
                           iterator_trap_0_port, QN => n271_port);
   iterator_trap_reg_29_inst : DFF_X1 port map( D => n410, CK => Clk, Q => 
                           iterator_trap_29_port, QN => n300);
   iterator_trap_reg_6_inst : DFF_X1 port map( D => n387, CK => Clk, Q => 
                           iterator_trap_6_port, QN => n277_port);
   iterator_trap_reg_17_inst : DFF_X1 port map( D => n398, CK => Clk, Q => 
                           iterator_trap_17_port, QN => n288);
   iterator_trap_reg_13_inst : DFF_X1 port map( D => n394, CK => Clk, Q => 
                           iterator_trap_13_port, QN => n284_port);
   iterator_trap_reg_9_inst : DFF_X1 port map( D => n390, CK => Clk, Q => 
                           iterator_trap_9_port, QN => n280_port);
   iterator_trap_reg_30_inst : DFF_X1 port map( D => n411, CK => Clk, Q => 
                           iterator_trap_30_port, QN => n301);
   iterator_trap_reg_26_inst : DFF_X1 port map( D => n407, CK => Clk, Q => 
                           iterator_trap_26_port, QN => n297);
   sig1_reg : DFF_X1 port map( D => n446, CK => Clk, Q => n188, QN => n517);
   s_trap_reg : DFF_X1 port map( D => n380, CK => Clk, Q => s_trap, QN => n339)
                           ;
   sig2_reg : DFF_X1 port map( D => n445, CK => Clk, Q => n140, QN => n_2379);
   iterator_ret_reg_0_inst : DFF_X1 port map( D => n413, CK => Clk, Q => 
                           iterator_ret_0_port, QN => n303);
   iterator_ret_reg_29_inst : DFF_X1 port map( D => n442, CK => Clk, Q => 
                           iterator_ret_29_port, QN => n332);
   iterator_ret_reg_27_inst : DFF_X1 port map( D => n440, CK => Clk, Q => 
                           iterator_ret_27_port, QN => n330);
   iterator_ret_reg_30_inst : DFF_X1 port map( D => n443, CK => Clk, Q => 
                           iterator_ret_30_port, QN => n333);
   iterator_ret_reg_22_inst : DFF_X1 port map( D => n435, CK => Clk, Q => 
                           iterator_ret_22_port, QN => n325);
   iterator_trap_reg_18_inst : DFF_X1 port map( D => n399, CK => Clk, Q => 
                           iterator_trap_18_port, QN => n289);
   iterator_trap_reg_14_inst : DFF_X1 port map( D => n395, CK => Clk, Q => 
                           iterator_trap_14_port, QN => n285);
   iterator_trap_reg_22_inst : DFF_X1 port map( D => n403, CK => Clk, Q => 
                           iterator_trap_22_port, QN => n293);
   iterator_trap_reg_21_inst : DFF_X1 port map( D => n402, CK => Clk, Q => 
                           iterator_trap_21_port, QN => n292);
   iterator_ret_reg_23_inst : DFF_X1 port map( D => n436, CK => Clk, Q => 
                           iterator_ret_23_port, QN => n326);
   iterator_ret_reg_18_inst : DFF_X1 port map( D => n431, CK => Clk, Q => 
                           iterator_ret_18_port, QN => n321);
   iterator_ret_reg_17_inst : DFF_X1 port map( D => n430, CK => Clk, Q => 
                           iterator_ret_17_port, QN => n320);
   iterator_ret_reg_15_inst : DFF_X1 port map( D => n428, CK => Clk, Q => 
                           iterator_ret_15_port, QN => n318);
   iterator_ret_reg_13_inst : DFF_X1 port map( D => n426, CK => Clk, Q => 
                           iterator_ret_13_port, QN => n316);
   iterator_ret_reg_12_inst : DFF_X1 port map( D => n425, CK => Clk, Q => 
                           iterator_ret_12_port, QN => n315);
   iterator_ret_reg_10_inst : DFF_X1 port map( D => n423, CK => Clk, Q => 
                           iterator_ret_10_port, QN => n313);
   iterator_ret_reg_9_inst : DFF_X1 port map( D => n422, CK => Clk, Q => 
                           iterator_ret_9_port, QN => n312);
   iterator_ret_reg_11_inst : DFF_X1 port map( D => n424, CK => Clk, Q => 
                           iterator_ret_11_port, QN => n314);
   iterator_trap_reg_4_inst : DFF_X1 port map( D => n385, CK => Clk, Q => 
                           iterator_trap_4_port, QN => n275_port);
   iterator_trap_reg_10_inst : DFF_X1 port map( D => n391, CK => Clk, Q => 
                           iterator_trap_10_port, QN => n281_port);
   iterator_trap_reg_27_inst : DFF_X1 port map( D => n408, CK => Clk, Q => 
                           iterator_trap_27_port, QN => n298);
   iterator_trap_reg_23_inst : DFF_X1 port map( D => n404, CK => Clk, Q => 
                           iterator_trap_23_port, QN => n294);
   iterator_trap_reg_20_inst : DFF_X1 port map( D => n401, CK => Clk, Q => 
                           iterator_trap_20_port, QN => n291);
   iterator_trap_reg_19_inst : DFF_X1 port map( D => n400, CK => Clk, Q => 
                           iterator_trap_19_port, QN => n290);
   iterator_ret_reg_2_inst : DFF_X1 port map( D => n415, CK => Clk, Q => 
                           iterator_ret_2_port, QN => n305);
   iterator_ret_reg_31_inst : DFF_X1 port map( D => n444, CK => Clk, Q => 
                           iterator_ret_31_port, QN => n334);
   iterator_ret_reg_6_inst : DFF_X1 port map( D => n419, CK => Clk, Q => 
                           iterator_ret_6_port, QN => n309);
   iterator_ret_reg_5_inst : DFF_X1 port map( D => n418, CK => Clk, Q => 
                           iterator_ret_5_port, QN => n308);
   iterator_ret_reg_4_inst : DFF_X1 port map( D => n417, CK => Clk, Q => 
                           iterator_ret_4_port, QN => n307);
   iterator_ret_reg_3_inst : DFF_X1 port map( D => n416, CK => Clk, Q => 
                           iterator_ret_3_port, QN => n306);
   iterator_ret_reg_1_inst : DFF_X1 port map( D => n414, CK => Clk, Q => 
                           iterator_ret_1_port, QN => n304);
   iterator_trap_reg_2_inst : DFF_X1 port map( D => n383, CK => Clk, Q => 
                           iterator_trap_2_port, QN => n273_port);
   iterator_trap_reg_1_inst : DFF_X1 port map( D => n382, CK => Clk, Q => 
                           iterator_trap_1_port, QN => n272_port);
   iterator_trap_reg_31_inst : DFF_X1 port map( D => n412, CK => Clk, Q => 
                           iterator_trap_31_port, QN => n302);
   iterator_trap_reg_7_inst : DFF_X1 port map( D => n388, CK => Clk, Q => 
                           iterator_trap_7_port, QN => n278_port);
   iterator_trap_reg_5_inst : DFF_X1 port map( D => n386, CK => Clk, Q => 
                           iterator_trap_5_port, QN => n276_port);
   iterator_trap_reg_3_inst : DFF_X1 port map( D => n384, CK => Clk, Q => 
                           iterator_trap_3_port, QN => n274_port);
   iterator_trap_reg_24_inst : DFF_X1 port map( D => n405, CK => Clk, Q => 
                           iterator_trap_24_port, QN => n295);
   iterator_trap_reg_16_inst : DFF_X1 port map( D => n397, CK => Clk, Q => 
                           iterator_trap_16_port, QN => n287);
   iterator_trap_reg_15_inst : DFF_X1 port map( D => n396, CK => Clk, Q => 
                           iterator_trap_15_port, QN => n286);
   iterator_trap_reg_12_inst : DFF_X1 port map( D => n393, CK => Clk, Q => 
                           iterator_trap_12_port, QN => n283_port);
   iterator_trap_reg_11_inst : DFF_X1 port map( D => n392, CK => Clk, Q => 
                           iterator_trap_11_port, QN => n282_port);
   iterator_trap_reg_8_inst : DFF_X1 port map( D => n389, CK => Clk, Q => 
                           iterator_trap_8_port, QN => n279_port);
   iterator_trap_reg_28_inst : DFF_X1 port map( D => n409, CK => Clk, Q => 
                           iterator_trap_28_port, QN => n299);
   iterator_trap_reg_25_inst : DFF_X1 port map( D => n406, CK => Clk, Q => 
                           iterator_trap_25_port, QN => n296);
   iterator_ret_reg_28_inst : DFF_X1 port map( D => n441, CK => Clk, Q => 
                           iterator_ret_28_port, QN => n331);
   iterator_ret_reg_25_inst : DFF_X1 port map( D => n438, CK => Clk, Q => 
                           iterator_ret_25_port, QN => n328);
   U3 : AND3_X2 port map( A1 => n27, A2 => n146_port, A3 => n147_port, ZN => 
                           n45_port);
   U4 : AND2_X2 port map( A1 => n152_port, A2 => n55_port, ZN => n1);
   U5 : INV_X1 port map( A => n1, ZN => n186);
   U6 : CLKBUF_X1 port map( A => N163, Z => n2);
   U7 : AND2_X1 port map( A1 => n196, A2 => n60_port, ZN => n31);
   U8 : AND2_X1 port map( A1 => n32, A2 => n194, ZN => n3);
   U9 : OR2_X1 port map( A1 => N54, A2 => N52, ZN => n4);
   U10 : BUF_X1 port map( A => n185, Z => n55_port);
   U11 : OR2_X1 port map( A1 => n199, A2 => n198, ZN => n5);
   U12 : INV_X1 port map( A => n31, ZN => n6);
   U13 : OR2_X1 port map( A1 => N162, A2 => N165, ZN => n7);
   U14 : CLKBUF_X1 port map( A => N175, Z => n8);
   U15 : INV_X1 port map( A => n26, ZN => n61_port);
   U16 : CLKBUF_X1 port map( A => N166, Z => n9);
   U17 : CLKBUF_X1 port map( A => N168, Z => n10);
   U18 : AND2_X1 port map( A1 => n33, A2 => n148_port, ZN => n11);
   U19 : CLKBUF_X1 port map( A => n38_port, Z => n12);
   U20 : CLKBUF_X1 port map( A => N57, Z => n13);
   U21 : OR2_X1 port map( A1 => N59, A2 => N58, ZN => n14);
   U22 : CLKBUF_X1 port map( A => N164, Z => n15);
   U23 : NAND2_X1 port map( A1 => n45_port, A2 => n11, ZN => n16);
   U24 : AND2_X1 port map( A1 => n17, A2 => n180, ZN => n146_port);
   U25 : NOR3_X1 port map( A1 => N173, A2 => N170, A3 => N171, ZN => n17);
   U26 : INV_X1 port map( A => N61, ZN => n18);
   U27 : BUF_X1 port map( A => n45_port, Z => n37_port);
   U28 : NOR3_X1 port map( A1 => N55, A2 => N53, A3 => n4, ZN => n190);
   U29 : NOR3_X1 port map( A1 => N164, A2 => N163, A3 => n7, ZN => n144);
   U30 : INV_X1 port map( A => n31, ZN => n19);
   U31 : INV_X1 port map( A => n31, ZN => n20);
   U32 : NOR3_X1 port map( A1 => n233, A2 => n230, A3 => n5, ZN => n195);
   U33 : AND2_X1 port map( A1 => n184, A2 => n46_port, ZN => n21);
   U34 : INV_X1 port map( A => n25, ZN => n22);
   U35 : INV_X1 port map( A => n25, ZN => n62_port);
   U36 : INV_X1 port map( A => n26, ZN => n23);
   U37 : NAND2_X1 port map( A1 => n140, A2 => n187, ZN => n24);
   U38 : NAND2_X1 port map( A1 => n24, A2 => n34_port, ZN => n445);
   U39 : AND2_X1 port map( A1 => n196, A2 => n60_port, ZN => n25);
   U40 : AND2_X1 port map( A1 => n196, A2 => n60_port, ZN => n26);
   U41 : AND2_X1 port map( A1 => n144, A2 => n145_port, ZN => n27);
   U42 : NOR3_X1 port map( A1 => N57, A2 => N56, A3 => n14, ZN => n191);
   U43 : NAND2_X1 port map( A1 => n45_port, A2 => n11, ZN => n184);
   U44 : INV_X1 port map( A => n26, ZN => n28);
   U45 : AND2_X1 port map( A1 => n16, A2 => n46_port, ZN => n151_port);
   U46 : NAND3_X1 port map( A1 => n21, A2 => n33, A3 => n37_port, ZN => n29);
   U47 : INV_X1 port map( A => n36_port, ZN => n30);
   U48 : BUF_X1 port map( A => n137, Z => n48_port);
   U49 : BUF_X1 port map( A => n137, Z => n47_port);
   U50 : BUF_X1 port map( A => n137, Z => n49_port);
   U51 : INV_X1 port map( A => n36_port, ZN => n56_port);
   U52 : BUF_X1 port map( A => n138, Z => n50_port);
   U53 : BUF_X1 port map( A => n138, Z => n51_port);
   U54 : BUF_X1 port map( A => n138, Z => n52_port);
   U55 : BUF_X1 port map( A => n238, Z => n58_port);
   U56 : BUF_X1 port map( A => n185, Z => n54_port);
   U57 : BUF_X1 port map( A => n185, Z => n53_port);
   U58 : BUF_X1 port map( A => n238, Z => n59_port);
   U59 : BUF_X1 port map( A => n238, Z => n60_port);
   U60 : AND2_X1 port map( A1 => n193, A2 => n192, ZN => n32);
   U61 : AND2_X1 port map( A1 => n143, A2 => n142, ZN => n33);
   U62 : BUF_X1 port map( A => Rst, Z => n64_port);
   U63 : BUF_X1 port map( A => Rst, Z => n63_port);
   U64 : BUF_X1 port map( A => Rst, Z => n65_port);
   U65 : INV_X1 port map( A => n39_port, ZN => n34_port);
   U66 : INV_X1 port map( A => n1, ZN => n35_port);
   U67 : AND2_X1 port map( A1 => n29, A2 => n55_port, ZN => n36_port);
   U68 : AND2_X1 port map( A1 => n29, A2 => n55_port, ZN => n39_port);
   U69 : INV_X1 port map( A => n12, ZN => n234);
   U70 : AND2_X1 port map( A1 => n191, A2 => n190, ZN => n38_port);
   U71 : NAND3_X1 port map( A1 => n195, A2 => n3, A3 => n38_port, ZN => n196);
   U72 : NAND4_X1 port map( A1 => n224, A2 => n225, A3 => n226, A4 => n223, ZN 
                           => n44_port);
   U73 : NOR3_X1 port map( A1 => n150_port, A2 => n149_port, A3 => N146, ZN => 
                           n46_port);
   U74 : INV_X1 port map( A => n39_port, ZN => n57_port);
   U75 : NAND2_X1 port map( A1 => IR_IN(26), A2 => IR_IN(27), ZN => n495);
   U76 : INV_X1 port map( A => n495, ZN => n241);
   U77 : INV_X1 port map( A => IR_IN(28), ZN => n244);
   U78 : INV_X1 port map( A => n491, ZN => n245);
   U79 : NAND3_X1 port map( A1 => n374, A2 => n244, A3 => n245, ZN => n246);
   U80 : NAND3_X1 port map( A1 => n457, A2 => n374, A3 => n244, ZN => n247);
   U81 : INV_X1 port map( A => IR_IN(31), ZN => n242);
   U82 : INV_X1 port map( A => IR_IN(30), ZN => n243);
   U83 : NAND4_X1 port map( A1 => IR_IN(29), A2 => IR_IN(28), A3 => n242, A4 =>
                           n243, ZN => n460);
   U84 : INV_X1 port map( A => n460, ZN => n240);
   U85 : NAND3_X1 port map( A1 => n65_port, A2 => n241, A3 => n240, ZN => n136)
                           ;
   U86 : INV_X1 port map( A => n136, ZN => n137);
   U87 : INV_X1 port map( A => N274, ZN => n116);
   U88 : INV_X1 port map( A => N273, ZN => n114);
   U89 : INV_X1 port map( A => N272, ZN => n112);
   U90 : INV_X1 port map( A => N271, ZN => n110);
   U91 : NAND4_X1 port map( A1 => n116, A2 => n114, A3 => n112, A4 => n110, ZN 
                           => n69);
   U92 : INV_X1 port map( A => N278, ZN => n124);
   U93 : INV_X1 port map( A => N277, ZN => n122);
   U94 : INV_X1 port map( A => N276, ZN => n120);
   U95 : INV_X1 port map( A => N275, ZN => n118);
   U96 : NAND4_X1 port map( A1 => n124, A2 => n122, A3 => n120, A4 => n118, ZN 
                           => n68);
   U97 : INV_X1 port map( A => N282, ZN => n132);
   U98 : INV_X1 port map( A => N281, ZN => n130);
   U99 : INV_X1 port map( A => N280, ZN => n128);
   U100 : INV_X1 port map( A => N279, ZN => n126);
   U101 : NAND4_X1 port map( A1 => n132, A2 => n130, A3 => n128, A4 => n126, ZN
                           => n67);
   U102 : INV_X1 port map( A => N284, ZN => n77);
   U103 : INV_X1 port map( A => N283, ZN => n134);
   U104 : NAND4_X1 port map( A1 => N254, A2 => N253, A3 => n77, A4 => n134, ZN 
                           => n66);
   U105 : NOR4_X1 port map( A1 => n69, A2 => n68, A3 => n67, A4 => n66, ZN => 
                           n75);
   U106 : INV_X1 port map( A => N258, ZN => n84);
   U107 : INV_X1 port map( A => N257, ZN => n82);
   U108 : INV_X1 port map( A => N256, ZN => n80);
   U109 : INV_X1 port map( A => N255, ZN => n79);
   U110 : NAND4_X1 port map( A1 => n84, A2 => n82, A3 => n80, A4 => n79, ZN => 
                           n73);
   U111 : INV_X1 port map( A => N262, ZN => n92);
   U112 : INV_X1 port map( A => N261, ZN => n90);
   U113 : INV_X1 port map( A => N260, ZN => n88);
   U114 : INV_X1 port map( A => N259, ZN => n86);
   U115 : NAND4_X1 port map( A1 => n92, A2 => n90, A3 => n88, A4 => n86, ZN => 
                           n72);
   U116 : INV_X1 port map( A => N266, ZN => n100);
   U117 : INV_X1 port map( A => N265, ZN => n98);
   U118 : INV_X1 port map( A => N264, ZN => n96);
   U119 : INV_X1 port map( A => N263, ZN => n94);
   U120 : NAND4_X1 port map( A1 => n100, A2 => n98, A3 => n96, A4 => n94, ZN =>
                           n71);
   U121 : INV_X1 port map( A => N270, ZN => n108);
   U122 : INV_X1 port map( A => N269, ZN => n106);
   U123 : INV_X1 port map( A => N268, ZN => n104);
   U124 : INV_X1 port map( A => N267, ZN => n102);
   U125 : NAND4_X1 port map( A1 => n108, A2 => n106, A3 => n104, A4 => n102, ZN
                           => n70);
   U126 : NOR4_X1 port map( A1 => n73, A2 => n72, A3 => n71, A4 => n70, ZN => 
                           n74);
   U127 : NAND2_X1 port map( A1 => n75, A2 => n74, ZN => n135);
   U128 : NAND2_X1 port map( A1 => n49_port, A2 => n135, ZN => n138);
   U129 : OAI22_X1 port map( A1 => n50_port, A2 => n77, B1 => n49_port, B2 => 
                           n76, ZN => n549);
   U130 : INV_X1 port map( A => N254, ZN => n78);
   U131 : OAI22_X1 port map( A1 => n78, A2 => n52_port, B1 => n49_port, B2 => 
                           n42_port, ZN => n548);
   U132 : OAI22_X1 port map( A1 => n50_port, A2 => n79, B1 => n49_port, B2 => 
                           n41_port, ZN => n547);
   U133 : OAI22_X1 port map( A1 => n51_port, A2 => n80, B1 => n49_port, B2 => 
                           n40_port, ZN => n546);
   U134 : OAI22_X1 port map( A1 => n51_port, A2 => n82, B1 => n49_port, B2 => 
                           n81, ZN => n545);
   U135 : OAI22_X1 port map( A1 => n50_port, A2 => n84, B1 => n49_port, B2 => 
                           n83, ZN => n544);
   U136 : OAI22_X1 port map( A1 => n51_port, A2 => n86, B1 => n49_port, B2 => 
                           n85, ZN => n543);
   U137 : OAI22_X1 port map( A1 => n50_port, A2 => n88, B1 => n49_port, B2 => 
                           n87, ZN => n542);
   U138 : OAI22_X1 port map( A1 => n50_port, A2 => n90, B1 => n48_port, B2 => 
                           n89, ZN => n541);
   U139 : OAI22_X1 port map( A1 => n50_port, A2 => n92, B1 => n48_port, B2 => 
                           n91, ZN => n540);
   U140 : OAI22_X1 port map( A1 => n50_port, A2 => n94, B1 => n48_port, B2 => 
                           n93, ZN => n539);
   U141 : OAI22_X1 port map( A1 => n51_port, A2 => n96, B1 => n48_port, B2 => 
                           n95, ZN => n538);
   U142 : OAI22_X1 port map( A1 => n50_port, A2 => n98, B1 => n48_port, B2 => 
                           n97, ZN => n537);
   U143 : OAI22_X1 port map( A1 => n51_port, A2 => n100, B1 => n48_port, B2 => 
                           n99, ZN => n536);
   U144 : OAI22_X1 port map( A1 => n50_port, A2 => n102, B1 => n48_port, B2 => 
                           n101, ZN => n535);
   U145 : OAI22_X1 port map( A1 => n51_port, A2 => n104, B1 => n48_port, B2 => 
                           n103, ZN => n534);
   U146 : OAI22_X1 port map( A1 => n51_port, A2 => n106, B1 => n48_port, B2 => 
                           n105, ZN => n533);
   U147 : OAI22_X1 port map( A1 => n50_port, A2 => n108, B1 => n48_port, B2 => 
                           n107, ZN => n532);
   U148 : OAI22_X1 port map( A1 => n51_port, A2 => n110, B1 => n48_port, B2 => 
                           n109, ZN => n531);
   U149 : OAI22_X1 port map( A1 => n52_port, A2 => n112, B1 => n48_port, B2 => 
                           n111, ZN => n530);
   U150 : OAI22_X1 port map( A1 => n52_port, A2 => n114, B1 => n47_port, B2 => 
                           n113, ZN => n529);
   U151 : OAI22_X1 port map( A1 => n52_port, A2 => n116, B1 => n47_port, B2 => 
                           n115, ZN => n528);
   U152 : OAI22_X1 port map( A1 => n52_port, A2 => n118, B1 => n47_port, B2 => 
                           n117, ZN => n527);
   U153 : OAI22_X1 port map( A1 => n50_port, A2 => n120, B1 => n47_port, B2 => 
                           n119, ZN => n526);
   U154 : OAI22_X1 port map( A1 => n52_port, A2 => n122, B1 => n47_port, B2 => 
                           n121, ZN => n525);
   U155 : OAI22_X1 port map( A1 => n52_port, A2 => n124, B1 => n47_port, B2 => 
                           n123, ZN => n524);
   U156 : OAI22_X1 port map( A1 => n52_port, A2 => n126, B1 => n47_port, B2 => 
                           n125, ZN => n523);
   U157 : OAI22_X1 port map( A1 => n52_port, A2 => n128, B1 => n47_port, B2 => 
                           n127, ZN => n522);
   U158 : OAI22_X1 port map( A1 => n51_port, A2 => n130, B1 => n47_port, B2 => 
                           n129, ZN => n521);
   U159 : OAI22_X1 port map( A1 => n51_port, A2 => n132, B1 => n47_port, B2 => 
                           n131, ZN => n520);
   U160 : OAI22_X1 port map( A1 => n51_port, A2 => n134, B1 => n47_port, B2 => 
                           n133, ZN => n519);
   U161 : OAI22_X1 port map( A1 => n136, A2 => n135, B1 => n336, B2 => n64_port
                           , ZN => n377);
   U162 : INV_X1 port map( A => N253, ZN => n139);
   U163 : OAI22_X1 port map( A1 => n139, A2 => n52_port, B1 => n47_port, B2 => 
                           n43_port, ZN => n518);
   U164 : INV_X1 port map( A => n247, ZN => n141);
   U165 : OAI21_X1 port map( B1 => n141, B2 => n140, A => n64_port, ZN => n187)
                           ;
   U166 : INV_X1 port map( A => n187, ZN => n185);
   U167 : INV_X1 port map( A => N153, ZN => n161_port);
   U168 : INV_X1 port map( A => N152, ZN => n160_port);
   U169 : INV_X1 port map( A => N151, ZN => n159_port);
   U170 : INV_X1 port map( A => N150, ZN => n158_port);
   U171 : NAND4_X1 port map( A1 => n161_port, A2 => n160_port, A3 => n159_port,
                           A4 => n158_port, ZN => n150_port);
   U172 : INV_X1 port map( A => N149, ZN => n157_port);
   U173 : INV_X1 port map( A => N148, ZN => n156_port);
   U174 : NAND2_X1 port map( A1 => n157_port, A2 => n156_port, ZN => n149_port)
                           ;
   U175 : NOR4_X1 port map( A1 => N160, A2 => N159, A3 => N158, A4 => N161, ZN 
                           => n143);
   U176 : NOR4_X1 port map( A1 => N154, A2 => N155, A3 => N156, A4 => N157, ZN 
                           => n142);
   U177 : NOR4_X1 port map( A1 => n150_port, A2 => n149_port, A3 => N145, A4 =>
                           N146, ZN => n148_port);
   U178 : INV_X1 port map( A => N147, ZN => n155_port);
   U179 : NOR4_X1 port map( A1 => N174, A2 => N175, A3 => N176, A4 => n155_port
                           , ZN => n147_port);
   U180 : NOR4_X1 port map( A1 => N168, A2 => N167, A3 => N166, A4 => N169, ZN 
                           => n145_port);
   U181 : NAND3_X1 port map( A1 => n151_port, A2 => n33, A3 => n37_port, ZN => 
                           n152_port);
   U182 : INV_X1 port map( A => N176, ZN => n153_port);
   U183 : OAI22_X1 port map( A1 => n56_port, A2 => n153_port, B1 => n334, B2 =>
                           n55_port, ZN => n444);
   U184 : INV_X1 port map( A => N146, ZN => n154_port);
   U185 : OAI22_X1 port map( A1 => n30, A2 => n154_port, B1 => n304, B2 => 
                           n55_port, ZN => n414);
   U186 : OAI22_X1 port map( A1 => n155_port, A2 => n57_port, B1 => n305, B2 =>
                           n55_port, ZN => n415);
   U187 : OAI22_X1 port map( A1 => n56_port, A2 => n156_port, B1 => n306, B2 =>
                           n55_port, ZN => n416);
   U188 : OAI22_X1 port map( A1 => n56_port, A2 => n157_port, B1 => n307, B2 =>
                           n55_port, ZN => n417);
   U189 : OAI22_X1 port map( A1 => n30, A2 => n158_port, B1 => n308, B2 => 
                           n55_port, ZN => n418);
   U190 : OAI22_X1 port map( A1 => n30, A2 => n159_port, B1 => n309, B2 => 
                           n55_port, ZN => n419);
   U191 : OAI22_X1 port map( A1 => n30, A2 => n160_port, B1 => n310, B2 => 
                           n54_port, ZN => n420);
   U192 : OAI22_X1 port map( A1 => n30, A2 => n161_port, B1 => n311, B2 => 
                           n54_port, ZN => n421);
   U193 : INV_X1 port map( A => N154, ZN => n162_port);
   U194 : OAI22_X1 port map( A1 => n35_port, A2 => n162_port, B1 => n312, B2 =>
                           n54_port, ZN => n422);
   U195 : INV_X1 port map( A => N155, ZN => n163_port);
   U196 : OAI22_X1 port map( A1 => n186, A2 => n163_port, B1 => n313, B2 => 
                           n54_port, ZN => n423);
   U197 : INV_X1 port map( A => N156, ZN => n164_port);
   U198 : OAI22_X1 port map( A1 => n35_port, A2 => n164_port, B1 => n314, B2 =>
                           n54_port, ZN => n424);
   U199 : INV_X1 port map( A => N157, ZN => n165_port);
   U200 : OAI22_X1 port map( A1 => n35_port, A2 => n165_port, B1 => n315, B2 =>
                           n54_port, ZN => n425);
   U201 : INV_X1 port map( A => N158, ZN => n166_port);
   U202 : OAI22_X1 port map( A1 => n186, A2 => n166_port, B1 => n316, B2 => 
                           n54_port, ZN => n426);
   U203 : INV_X1 port map( A => N159, ZN => n167_port);
   U204 : OAI22_X1 port map( A1 => n56_port, A2 => n167_port, B1 => n317, B2 =>
                           n54_port, ZN => n427);
   U205 : INV_X1 port map( A => N160, ZN => n168_port);
   U206 : OAI22_X1 port map( A1 => n35_port, A2 => n168_port, B1 => n318, B2 =>
                           n54_port, ZN => n428);
   U207 : INV_X1 port map( A => N161, ZN => n169_port);
   U208 : OAI22_X1 port map( A1 => n34_port, A2 => n169_port, B1 => n319, B2 =>
                           n54_port, ZN => n429);
   U209 : INV_X1 port map( A => N162, ZN => n170_port);
   U210 : OAI22_X1 port map( A1 => n35_port, A2 => n170_port, B1 => n320, B2 =>
                           n54_port, ZN => n430);
   U211 : INV_X1 port map( A => n2, ZN => n171_port);
   U212 : OAI22_X1 port map( A1 => n186, A2 => n171_port, B1 => n321, B2 => 
                           n53_port, ZN => n431);
   U213 : INV_X1 port map( A => n15, ZN => n172_port);
   U214 : OAI22_X1 port map( A1 => n34_port, A2 => n172_port, B1 => n322, B2 =>
                           n53_port, ZN => n432);
   U215 : INV_X1 port map( A => N165, ZN => n173_port);
   U216 : OAI22_X1 port map( A1 => n56_port, A2 => n173_port, B1 => n323, B2 =>
                           n53_port, ZN => n433);
   U217 : INV_X1 port map( A => n9, ZN => n174_port);
   U218 : OAI22_X1 port map( A1 => n34_port, A2 => n174_port, B1 => n324, B2 =>
                           n53_port, ZN => n434);
   U219 : INV_X1 port map( A => N167, ZN => n175_port);
   U220 : OAI22_X1 port map( A1 => n57_port, A2 => n175_port, B1 => n325, B2 =>
                           n53_port, ZN => n435);
   U221 : INV_X1 port map( A => n10, ZN => n176_port);
   U222 : OAI22_X1 port map( A1 => n186, A2 => n176_port, B1 => n326, B2 => 
                           n54_port, ZN => n436);
   U223 : INV_X1 port map( A => N169, ZN => n177);
   U224 : OAI22_X1 port map( A1 => n56_port, A2 => n177, B1 => n327, B2 => 
                           n53_port, ZN => n437);
   U225 : INV_X1 port map( A => N170, ZN => n178);
   U226 : OAI22_X1 port map( A1 => n34_port, A2 => n178, B1 => n328, B2 => 
                           n53_port, ZN => n438);
   U227 : INV_X1 port map( A => N171, ZN => n179);
   U228 : OAI22_X1 port map( A1 => n30, A2 => n179, B1 => n329, B2 => n53_port,
                           ZN => n439);
   U229 : INV_X1 port map( A => N172, ZN => n180);
   U230 : OAI22_X1 port map( A1 => n57_port, A2 => n180, B1 => n330, B2 => 
                           n53_port, ZN => n440);
   U231 : INV_X1 port map( A => N173, ZN => n181);
   U232 : OAI22_X1 port map( A1 => n34_port, A2 => n181, B1 => n331, B2 => 
                           n53_port, ZN => n441);
   U233 : INV_X1 port map( A => N174, ZN => n182);
   U234 : OAI22_X1 port map( A1 => n57_port, A2 => n182, B1 => n332, B2 => 
                           n53_port, ZN => n442);
   U235 : INV_X1 port map( A => n8, ZN => n183);
   U236 : OAI22_X1 port map( A1 => n57_port, A2 => n183, B1 => n333, B2 => 
                           n53_port, ZN => n443);
   U237 : OAI22_X1 port map( A1 => n187, A2 => n16, B1 => n340, B2 => n64_port,
                           ZN => n379);
   U238 : MUX2_X1 port map( A => n187, B => n1, S => n303, Z => n413);
   U239 : INV_X1 port map( A => n246, ZN => n189);
   U240 : OAI21_X1 port map( B1 => n189, B2 => n188, A => n64_port, ZN => n239)
                           ;
   U241 : INV_X1 port map( A => n239, ZN => n238);
   U242 : INV_X1 port map( A => N63, ZN => n226);
   U243 : INV_X1 port map( A => N62, ZN => n225);
   U244 : INV_X1 port map( A => N61, ZN => n224);
   U245 : INV_X1 port map( A => N60, ZN => n223);
   U246 : NAND4_X1 port map( A1 => n226, A2 => n225, A3 => n18, A4 => n223, ZN 
                           => n233);
   U247 : INV_X1 port map( A => N65, ZN => n197);
   U248 : INV_X1 port map( A => N64, ZN => n227);
   U249 : NAND2_X1 port map( A1 => n197, A2 => n227, ZN => n230);
   U250 : INV_X1 port map( A => N35, ZN => n198);
   U251 : INV_X1 port map( A => N36, ZN => n199);
   U252 : NOR4_X1 port map( A1 => N51, A2 => N49, A3 => N50, A4 => N48, ZN => 
                           n193);
   U253 : NOR4_X1 port map( A1 => N44, A2 => N45, A3 => N46, A4 => N47, ZN => 
                           n192);
   U254 : INV_X1 port map( A => N43, ZN => n206);
   U255 : INV_X1 port map( A => N42, ZN => n205);
   U256 : INV_X1 port map( A => N41, ZN => n204);
   U257 : INV_X1 port map( A => N40, ZN => n203);
   U258 : NAND4_X1 port map( A1 => n206, A2 => n205, A3 => n204, A4 => n203, ZN
                           => n229);
   U259 : INV_X1 port map( A => N39, ZN => n202);
   U260 : INV_X1 port map( A => N38, ZN => n201);
   U261 : NAND2_X1 port map( A1 => n202, A2 => n201, ZN => n228);
   U262 : NOR4_X1 port map( A1 => n229, A2 => n228, A3 => N34, A4 => N37, ZN =>
                           n194);
   U263 : OAI22_X1 port map( A1 => n61_port, A2 => n197, B1 => n302, B2 => 
                           n60_port, ZN => n412);
   U264 : OAI22_X1 port map( A1 => n198, A2 => n20, B1 => n272_port, B2 => 
                           n60_port, ZN => n382);
   U265 : OAI22_X1 port map( A1 => n199, A2 => n6, B1 => n273_port, B2 => 
                           n60_port, ZN => n383);
   U266 : INV_X1 port map( A => N37, ZN => n200);
   U267 : OAI22_X1 port map( A1 => n23, A2 => n200, B1 => n274_port, B2 => 
                           n60_port, ZN => n384);
   U268 : OAI22_X1 port map( A1 => n20, A2 => n201, B1 => n275_port, B2 => 
                           n60_port, ZN => n385);
   U269 : OAI22_X1 port map( A1 => n61_port, A2 => n202, B1 => n276_port, B2 =>
                           n60_port, ZN => n386);
   U270 : OAI22_X1 port map( A1 => n22, A2 => n203, B1 => n277_port, B2 => 
                           n60_port, ZN => n387);
   U271 : OAI22_X1 port map( A1 => n23, A2 => n204, B1 => n278_port, B2 => 
                           n60_port, ZN => n388);
   U272 : OAI22_X1 port map( A1 => n61_port, A2 => n205, B1 => n279_port, B2 =>
                           n59_port, ZN => n389);
   U273 : OAI22_X1 port map( A1 => n62_port, A2 => n206, B1 => n280_port, B2 =>
                           n59_port, ZN => n390);
   U274 : INV_X1 port map( A => N44, ZN => n207);
   U275 : OAI22_X1 port map( A1 => n19, A2 => n207, B1 => n281_port, B2 => 
                           n59_port, ZN => n391);
   U276 : INV_X1 port map( A => N45, ZN => n208);
   U277 : OAI22_X1 port map( A1 => n28, A2 => n208, B1 => n282_port, B2 => 
                           n59_port, ZN => n392);
   U278 : INV_X1 port map( A => N46, ZN => n209);
   U279 : OAI22_X1 port map( A1 => n23, A2 => n209, B1 => n283_port, B2 => 
                           n59_port, ZN => n393);
   U280 : INV_X1 port map( A => N47, ZN => n210);
   U281 : OAI22_X1 port map( A1 => n22, A2 => n210, B1 => n284_port, B2 => 
                           n59_port, ZN => n394);
   U282 : INV_X1 port map( A => N48, ZN => n211);
   U283 : OAI22_X1 port map( A1 => n62_port, A2 => n211, B1 => n285, B2 => 
                           n59_port, ZN => n395);
   U284 : INV_X1 port map( A => N49, ZN => n212);
   U285 : OAI22_X1 port map( A1 => n28, A2 => n212, B1 => n286, B2 => n59_port,
                           ZN => n396);
   U286 : INV_X1 port map( A => N50, ZN => n213);
   U287 : OAI22_X1 port map( A1 => n61_port, A2 => n213, B1 => n287, B2 => 
                           n59_port, ZN => n397);
   U288 : INV_X1 port map( A => N51, ZN => n214);
   U289 : OAI22_X1 port map( A1 => n22, A2 => n214, B1 => n288, B2 => n59_port,
                           ZN => n398);
   U290 : INV_X1 port map( A => N52, ZN => n215);
   U291 : OAI22_X1 port map( A1 => n6, A2 => n215, B1 => n289, B2 => n59_port, 
                           ZN => n399);
   U292 : INV_X1 port map( A => N53, ZN => n216);
   U293 : OAI22_X1 port map( A1 => n20, A2 => n216, B1 => n290, B2 => n58_port,
                           ZN => n400);
   U294 : INV_X1 port map( A => N54, ZN => n217);
   U295 : OAI22_X1 port map( A1 => n19, A2 => n217, B1 => n291, B2 => n58_port,
                           ZN => n401);
   U296 : INV_X1 port map( A => N55, ZN => n218);
   U297 : OAI22_X1 port map( A1 => n22, A2 => n218, B1 => n292, B2 => n58_port,
                           ZN => n402);
   U298 : INV_X1 port map( A => N56, ZN => n219);
   U299 : OAI22_X1 port map( A1 => n19, A2 => n219, B1 => n293, B2 => n58_port,
                           ZN => n403);
   U300 : INV_X1 port map( A => n13, ZN => n220);
   U301 : OAI22_X1 port map( A1 => n19, A2 => n220, B1 => n294, B2 => n58_port,
                           ZN => n404);
   U302 : INV_X1 port map( A => N58, ZN => n221);
   U303 : OAI22_X1 port map( A1 => n28, A2 => n221, B1 => n295, B2 => n59_port,
                           ZN => n405);
   U304 : INV_X1 port map( A => N59, ZN => n222);
   U305 : OAI22_X1 port map( A1 => n23, A2 => n222, B1 => n296, B2 => n58_port,
                           ZN => n406);
   U306 : OAI22_X1 port map( A1 => n62_port, A2 => n223, B1 => n297, B2 => 
                           n58_port, ZN => n407);
   U307 : OAI22_X1 port map( A1 => n20, A2 => n224, B1 => n298, B2 => n58_port,
                           ZN => n408);
   U308 : OAI22_X1 port map( A1 => n28, A2 => n225, B1 => n299, B2 => n58_port,
                           ZN => n409);
   U309 : OAI22_X1 port map( A1 => n6, A2 => n226, B1 => n300, B2 => n58_port, 
                           ZN => n410);
   U310 : OAI22_X1 port map( A1 => n62_port, A2 => n227, B1 => n301, B2 => 
                           n58_port, ZN => n411);
   U311 : NOR4_X1 port map( A1 => n229, A2 => n228, A3 => N37, A4 => N35, ZN =>
                           n236);
   U312 : INV_X1 port map( A => n230, ZN => n231);
   U313 : NAND4_X1 port map( A1 => N34, A2 => N36, A3 => n58_port, A4 => n231, 
                           ZN => n232);
   U314 : NOR3_X1 port map( A1 => n234, A2 => n44_port, A3 => n232, ZN => n235)
                           ;
   U315 : NAND3_X1 port map( A1 => n236, A2 => n32, A3 => n235, ZN => n237);
   U316 : OAI21_X1 port map( B1 => n339, B2 => n65_port, A => n237, ZN => n380)
                           ;
   U317 : OAI21_X1 port map( B1 => n517, B2 => n60_port, A => n6, ZN => n446);
   U318 : MUX2_X1 port map( A => n239, B => n25, S => n271_port, Z => n381);
   U319 : MUX2_X1 port map( A => sb_op_port, B => n248, S => n63_port, Z => 
                           n345);
   U320 : MUX2_X1 port map( A => n249, B => signed_unsigned_i, S => n63_port, Z
                           => n344);
   U321 : MUX2_X1 port map( A => signed_unsigned_port, B => n249, S => n63_port
                           , Z => n343);
   U322 : INV_X1 port map( A => n250, ZN => aluOpcode_i_5_port);
   U323 : AOI211_X1 port map( C1 => n241, C2 => n251, A => n252, B => n253_port
                           , ZN => n250);
   U324 : OAI211_X1 port map( C1 => n254_port, C2 => n255_port, A => n246, B =>
                           n247, ZN => n253_port);
   U325 : AND4_X1 port map( A1 => n256_port, A2 => n257_port, A3 => n258_port, 
                           A4 => n259_port, ZN => n255_port);
   U326 : OR2_X1 port map( A1 => n260_port, A2 => n261_port, ZN => n257_port);
   U327 : NAND4_X1 port map( A1 => n246, A2 => n262_port, A3 => n247, A4 => 
                           n263_port, ZN => aluOpcode_i_4_port);
   U328 : AOI211_X1 port map( C1 => n264_port, C2 => n265_port, A => n266_port,
                           B => n267_port, ZN => n263_port);
   U329 : INV_X1 port map( A => n268_port, ZN => n267_port);
   U330 : OAI21_X1 port map( B1 => n269_port, B2 => n270_port, A => n335, ZN =>
                           n265_port);
   U331 : NAND4_X1 port map( A1 => n337, A2 => n338, A3 => n341, A4 => n342, ZN
                           => aluOpcode_i_3_port);
   U332 : AOI211_X1 port map( C1 => n264_port, C2 => n346, A => n347, B => n348
                           , ZN => n342);
   U333 : OAI221_X1 port map( B1 => n349, B2 => n269_port, C1 => n350, C2 => 
                           n351, A => n335, ZN => n346);
   U334 : NAND4_X1 port map( A1 => n352, A2 => n353, A3 => n354, A4 => n355, ZN
                           => aluOpcode_i_2_port);
   U335 : AOI211_X1 port map( C1 => n356, C2 => n245, A => n357, B => n358, ZN 
                           => n355);
   U336 : INV_X1 port map( A => n359, ZN => n358);
   U337 : AOI21_X1 port map( B1 => n264_port, B2 => n360, A => n361, ZN => n354
                           );
   U338 : OAI221_X1 port map( B1 => n261_port, B2 => n362, C1 => n363, C2 => 
                           n349, A => n364, ZN => n360);
   U339 : NAND4_X1 port map( A1 => n365, A2 => n337, A3 => n366, A4 => n367, ZN
                           => aluOpcode_i_1_port);
   U340 : AOI221_X1 port map( B1 => n264_port, B2 => n368, C1 => n251, C2 => 
                           n369, A => n370, ZN => n367);
   U341 : NAND3_X1 port map( A1 => n246, A2 => n352, A3 => n371, ZN => n370);
   U342 : INV_X1 port map( A => n248, ZN => n371);
   U343 : NAND3_X1 port map( A1 => n372, A2 => n264_port, A3 => n373, ZN => 
                           n352);
   U344 : INV_X1 port map( A => n375, ZN => n369);
   U345 : OAI21_X1 port map( B1 => n363, B2 => n260_port, A => n376, ZN => n368
                           );
   U346 : AOI22_X1 port map( A1 => n378, A2 => n245, B1 => n447, B2 => n241, ZN
                           => n366);
   U347 : AOI22_X1 port map( A1 => n448, A2 => n264_port, B1 => n449, B2 => 
                           n356, ZN => n337);
   U348 : INV_X1 port map( A => n450, ZN => n365);
   U349 : NAND4_X1 port map( A1 => n451, A2 => n452, A3 => n453, A4 => n454, ZN
                           => aluOpcode_i_0_port);
   U350 : AOI221_X1 port map( B1 => n251, B2 => n449, C1 => n455, C2 => n245, A
                           => n450, ZN => n454);
   U351 : NAND4_X1 port map( A1 => n341, A2 => n247, A3 => n456, A4 => n353, ZN
                           => n450);
   U352 : AOI21_X1 port map( B1 => n264_port, B2 => n458, A => n459, ZN => n453
                           );
   U353 : AOI21_X1 port map( B1 => n460, B2 => n461, A => n462, ZN => n459);
   U354 : NAND4_X1 port map( A1 => n256_port, A2 => n463, A3 => n464, A4 => 
                           n465, ZN => n458);
   U355 : AOI21_X1 port map( B1 => n466, B2 => n467, A => n468, ZN => n465);
   U356 : INV_X1 port map( A => n469, ZN => n464);
   U357 : AOI21_X1 port map( B1 => n470, B2 => n349, A => n269_port, ZN => n469
                           );
   U358 : INV_X1 port map( A => n467, ZN => n349);
   U359 : NAND2_X1 port map( A1 => n270_port, A2 => n260_port, ZN => n467);
   U360 : NAND3_X1 port map( A1 => IR_IN(31), A2 => IR_IN(30), A3 => n471, ZN 
                           => n452);
   U361 : OAI21_X1 port map( B1 => n378, B2 => n356, A => n457, ZN => n451);
   U362 : NAND4_X1 port map( A1 => n341, A2 => n472, A3 => n473, A4 => 
                           n262_port, ZN => N551);
   U363 : OAI211_X1 port map( C1 => n474, C2 => n475, A => n244, B => n476, ZN 
                           => n473);
   U364 : NOR2_X1 port map( A1 => n477, A2 => n462, ZN => n475);
   U365 : NOR4_X1 port map( A1 => IR_IN(31), A2 => IR_IN(30), A3 => n478, A4 =>
                           n479, ZN => n474);
   U366 : AOI21_X1 port map( B1 => n480, B2 => n481, A => n482, ZN => n478);
   U367 : INV_X1 port map( A => n266_port, ZN => n472);
   U368 : AOI21_X1 port map( B1 => n240, B2 => n457, A => n361, ZN => n341);
   U369 : NAND4_X1 port map( A1 => n483, A2 => n484, A3 => n485, A4 => n486, ZN
                           => N550);
   U370 : NOR3_X1 port map( A1 => n487, A2 => n266_port, A3 => n357, ZN => n486
                           );
   U371 : OAI211_X1 port map( C1 => n460, C2 => n479, A => n268_port, B => n488
                           , ZN => n357);
   U372 : AOI221_X1 port map( B1 => n251, B2 => n241, C1 => n356, C2 => n489, A
                           => n348, ZN => n488);
   U373 : AOI22_X1 port map( A1 => n245, A2 => n447, B1 => n490, B2 => n378, ZN
                           => n268_port);
   U374 : NOR3_X1 port map( A1 => n476, A2 => n244, A3 => n477, ZN => n378);
   U375 : OAI211_X1 port map( C1 => n460, C2 => n491, A => n338, B => n492, ZN 
                           => n266_port);
   U376 : AOI221_X1 port map( B1 => n251, B2 => n457, C1 => n489, C2 => n487, A
                           => n493, ZN => n492);
   U377 : INV_X1 port map( A => n353, ZN => n493);
   U378 : NAND3_X1 port map( A1 => IR_IN(31), A2 => n241, A3 => n494, ZN => 
                           n353);
   U379 : INV_X1 port map( A => n496, ZN => n251);
   U395 : AOI21_X1 port map( B1 => n245, B2 => n356, A => n497, ZN => n338);
   U396 : NOR3_X1 port map( A1 => n495, A2 => IR_IN(30), A3 => n498, ZN => n497
                           );
   U397 : NAND2_X1 port map( A1 => n460, A2 => n496, ZN => n487);
   U398 : NAND2_X1 port map( A1 => n374, A2 => IR_IN(28), ZN => n496);
   U399 : NOR2_X1 port map( A1 => n477, A2 => IR_IN(29), ZN => n374);
   U400 : AOI21_X1 port map( B1 => n264_port, B2 => n499, A => n252, ZN => n485
                           );
   U401 : OR3_X1 port map( A1 => n361, A2 => n500, A3 => n347, ZN => n252);
   U402 : OAI211_X1 port map( C1 => n375, C2 => n461, A => n456, B => n359, ZN 
                           => n347);
   U403 : AOI21_X1 port map( B1 => IR_IN(31), B2 => n348, A => n248, ZN => n359
                           );
   U404 : NOR4_X1 port map( A1 => n242, A2 => n498, A3 => n479, A4 => IR_IN(30)
                           , ZN => n248);
   U405 : AND2_X1 port map( A1 => n455, A2 => n490, ZN => n348);
   U406 : NAND2_X1 port map( A1 => n479, A2 => n491, ZN => n490);
   U407 : INV_X1 port map( A => n457, ZN => n479);
   U408 : NOR3_X1 port map( A1 => IR_IN(29), A2 => IR_IN(30), A3 => n244, ZN =>
                           n455);
   U409 : NAND3_X1 port map( A1 => IR_IN(31), A2 => n457, A3 => n494, ZN => 
                           n456);
   U410 : INV_X1 port map( A => n447, ZN => n461);
   U411 : NOR2_X1 port map( A1 => n498, A2 => n477, ZN => n447);
   U412 : NAND2_X1 port map( A1 => IR_IN(30), A2 => n242, ZN => n477);
   U413 : NOR2_X1 port map( A1 => n449, A2 => n457, ZN => n375);
   U414 : INV_X1 port map( A => n262_port, ZN => n500);
   U415 : OAI211_X1 port map( C1 => n501, C2 => n471, A => IR_IN(30), B => 
                           IR_IN(31), ZN => n262_port);
   U416 : NOR3_X1 port map( A1 => n476, A2 => n244, A3 => n491, ZN => n471);
   U417 : NAND2_X1 port map( A1 => IR_IN(26), A2 => n502, ZN => n491);
   U418 : INV_X1 port map( A => IR_IN(29), ZN => n476);
   U419 : NOR2_X1 port map( A1 => n495, A2 => n498, ZN => n501);
   U420 : NOR4_X1 port map( A1 => n462, A2 => n242, A3 => n498, A4 => n243, ZN 
                           => n361);
   U421 : NAND4_X1 port map( A1 => n260_port, A2 => n270_port, A3 => n335, A4 
                           => n503, ZN => n499);
   U422 : NOR2_X1 port map( A1 => n482, A2 => n448, ZN => n503);
   U423 : OAI22_X1 port map( A1 => n269_port, A2 => n470, B1 => n470, B2 => 
                           n504, ZN => n448);
   U424 : NAND3_X1 port map( A1 => n505, A2 => n506, A3 => IR_IN(2), ZN => n470
                           );
   U425 : INV_X1 port map( A => n507, ZN => n269_port);
   U426 : OAI211_X1 port map( C1 => n363, C2 => n351, A => n256_port, B => n376
                           , ZN => n482);
   U427 : AOI211_X1 port map( C1 => n507, C2 => n480, A => n468, B => n508, ZN 
                           => n376);
   U428 : OAI21_X1 port map( B1 => n362, B2 => n504, A => n258_port, ZN => n508
                           );
   U429 : NAND4_X1 port map( A1 => n481, A2 => IR_IN(4), A3 => n505, A4 => n509
                           , ZN => n258_port);
   U430 : INV_X1 port map( A => n372, ZN => n504);
   U431 : OAI211_X1 port map( C1 => n350, C2 => n362, A => n364, B => n259_port
                           , ZN => n468);
   U432 : NAND4_X1 port map( A1 => IR_IN(4), A2 => IR_IN(2), A3 => n507, A4 => 
                           n505, ZN => n259_port);
   U433 : NAND2_X1 port map( A1 => n373, A2 => n507, ZN => n364);
   U434 : INV_X1 port map( A => n351, ZN => n373);
   U435 : INV_X1 port map( A => n510, ZN => n362);
   U436 : NOR2_X1 port map( A1 => n511, A2 => IR_IN(1), ZN => n507);
   U437 : NAND4_X1 port map( A1 => n466, A2 => IR_IN(4), A3 => n505, A4 => n509
                           , ZN => n256_port);
   U438 : NAND2_X1 port map( A1 => n512, A2 => IR_IN(2), ZN => n351);
   U439 : INV_X1 port map( A => n513, ZN => n335);
   U440 : OAI21_X1 port map( B1 => n363, B2 => n260_port, A => n463, ZN => n513
                           );
   U441 : OAI21_X1 port map( B1 => n480, B2 => n510, A => n481, ZN => n463);
   U442 : INV_X1 port map( A => n261_port, ZN => n481);
   U443 : NAND2_X1 port map( A1 => IR_IN(1), A2 => IR_IN(0), ZN => n261_port);
   U444 : NOR4_X1 port map( A1 => n509, A2 => IR_IN(3), A3 => IR_IN(4), A4 => 
                           IR_IN(5), ZN => n510);
   U445 : INV_X1 port map( A => n270_port, ZN => n480);
   U446 : NOR2_X1 port map( A1 => n466, A2 => n372, ZN => n363);
   U447 : NOR2_X1 port map( A1 => IR_IN(0), A2 => IR_IN(1), ZN => n372);
   U448 : INV_X1 port map( A => n350, ZN => n466);
   U449 : NAND2_X1 port map( A1 => IR_IN(1), A2 => n511, ZN => n350);
   U450 : INV_X1 port map( A => IR_IN(0), ZN => n511);
   U451 : NAND2_X1 port map( A1 => n512, A2 => n509, ZN => n270_port);
   U452 : NOR3_X1 port map( A1 => IR_IN(3), A2 => IR_IN(4), A3 => n514, ZN => 
                           n512);
   U453 : INV_X1 port map( A => IR_IN(5), ZN => n514);
   U454 : NAND3_X1 port map( A1 => n509, A2 => n506, A3 => n505, ZN => 
                           n260_port);
   U455 : AND2_X1 port map( A1 => IR_IN(5), A2 => IR_IN(3), ZN => n505);
   U456 : INV_X1 port map( A => IR_IN(4), ZN => n506);
   U457 : INV_X1 port map( A => IR_IN(2), ZN => n509);
   U458 : INV_X1 port map( A => n254_port, ZN => n264_port);
   U459 : NAND4_X1 port map( A1 => n494, A2 => n457, A3 => n515, A4 => n516, ZN
                           => n254_port);
   U460 : NOR4_X1 port map( A1 => IR_IN(31), A2 => IR_IN(9), A3 => IR_IN(8), A4
                           => IR_IN(7), ZN => n516);
   U461 : NOR2_X1 port map( A1 => IR_IN(6), A2 => IR_IN(10), ZN => n515);
   U462 : NOR2_X1 port map( A1 => IR_IN(26), A2 => IR_IN(27), ZN => n457);
   U463 : NOR3_X1 port map( A1 => IR_IN(29), A2 => IR_IN(30), A3 => IR_IN(28), 
                           ZN => n494);
   U464 : INV_X1 port map( A => n356, ZN => n484);
   U465 : NOR3_X1 port map( A1 => IR_IN(30), A2 => IR_IN(31), A3 => n498, ZN =>
                           n356);
   U466 : NAND2_X1 port map( A1 => IR_IN(29), A2 => n244, ZN => n498);
   U467 : NAND3_X1 port map( A1 => n244, A2 => n242, A3 => n449, ZN => n483);
   U468 : NAND2_X1 port map( A1 => n462, A2 => n495, ZN => n449);
   U469 : INV_X1 port map( A => n489, ZN => n462);
   U470 : NOR2_X1 port map( A1 => n502, A2 => IR_IN(26), ZN => n489);
   U471 : INV_X1 port map( A => IR_IN(27), ZN => n502);

end SYN_dlx_cu_hw;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity DLX_IR_SIZE32_PC_SIZE32 is

   port( CLK, RST : in std_logic;  IRAM_ADDRESS : out std_logic_vector (31 
         downto 0);  IRAM_ISSUE : out std_logic;  IRAM_READY : in std_logic;  
         IRAM_DATA : in std_logic_vector (63 downto 0);  DRAM_ADDRESS : out 
         std_logic_vector (31 downto 0);  DRAM_ISSUE, DRAM_READNOTWRITE : out 
         std_logic;  DRAM_READY : in std_logic;  DRAM_DATA : inout 
         std_logic_vector (63 downto 0));

end DLX_IR_SIZE32_PC_SIZE32;

architecture SYN_dlx_rtl of DLX_IR_SIZE32_PC_SIZE32 is

   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component TBUF_X1
      port( A, EN : in std_logic;  Z : out std_logic);
   end component;
   
   component DATAPTH_NBIT32_REG_BIT5
      port( CLK, RST : in std_logic;  PC, IR : in std_logic_vector (31 downto 
            0);  PC_OUT : out std_logic_vector (31 downto 0);  NPC_LATCH_EN, 
            ir_LATCH_EN, signed_op, trap_cs, ret_cs, RF1, RF2, WF1, 
            regImm_LATCH_EN, S1, S2, EN2, lhi_sel, jump_en, branch_cond, sb_op,
            RM, WM, EN3, S3 : in std_logic;  instruction_alu : in 
            std_logic_vector (0 to 5);  DATA_MEM_ADDR, DATA_MEM_IN : out 
            std_logic_vector (31 downto 0);  DATA_MEM_OUT : in std_logic_vector
            (31 downto 0);  DATA_MEM_ENABLE, DATA_MEM_RM, DATA_MEM_WM : out 
            std_logic);
   end component;
   
   component 
      dlx_cu_MICROCODE_MEM_SIZE62_FUNC_SIZE11_OP_CODE_SIZE6_IR_SIZE32_CW_SIZE15
      port( Clk, Rst : in std_logic;  IR_IN : in std_logic_vector (31 downto 0)
            ;  IR_LATCH_EN, NPC_LATCH_EN, RegA_LATCH_EN, RegB_LATCH_EN, 
            RegIMM_LATCH_EN, MUXA_SEL, MUXB_SEL, ALU_OUTREG_EN, EQ_COND : out 
            std_logic;  ALU_OPCODE : out std_logic_vector (0 to 5);  
            signed_unsigned, DRAM_WE, LMD_LATCH_EN, JUMP_EN, PC_LATCH_EN, 
            WB_MUX_SEL, RF_WE, lhi_sel, sb_op, s_trap, s_ret : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal IR_31_port, IR_30_port, IR_29_port, IR_28_port, IR_27_port, 
      IR_26_port, IR_25_port, IR_24_port, IR_23_port, IR_22_port, IR_21_port, 
      IR_20_port, IR_19_port, IR_18_port, IR_17_port, IR_16_port, IR_15_port, 
      IR_14_port, IR_13_port, IR_12_port, IR_11_port, IR_10_port, IR_9_port, 
      IR_8_port, IR_7_port, IR_6_port, IR_5_port, IR_4_port, IR_3_port, 
      IR_2_port, IR_1_port, IR_0_port, IR_LATCH_EN_i, PC_31_port, PC_30_port, 
      PC_29_port, PC_28_port, PC_27_port, PC_26_port, PC_25_port, PC_24_port, 
      PC_23_port, PC_22_port, PC_21_port, PC_20_port, PC_19_port, PC_18_port, 
      PC_17_port, PC_16_port, PC_15_port, PC_14_port, PC_13_port, PC_12_port, 
      PC_11_port, PC_10_port, PC_9_port, PC_8_port, PC_7_port, PC_6_port, 
      PC_5_port, PC_4_port, PC_3_port, PC_2_port, PC_1_port, PC_0_port, 
      PC_LATCH_EN_i, NPC_LATCH_EN_i, RegA_LATCH_EN_i, RegB_LATCH_EN_i, 
      RegIMM_LATCH_EN_i, MUXA_SEL_i, MUXB_SEL_i, ALU_OUTREG_EN_i, EQ_COND_i, 
      ALU_OPCODE_i_5_port, ALU_OPCODE_i_4_port, ALU_OPCODE_i_3_port, 
      ALU_OPCODE_i_2_port, ALU_OPCODE_i_1_port, ALU_OPCODE_i_0_port, 
      signed_unsigned_i, DRAM_WE_i, LMD_LATCH_EN_i, JUMP_EN_i, WB_MUX_SEL_i, 
      RF_WE_i, lhi_sel_i, sb_op_i, trap_cs_i, ret_cs_i, DATA_MEM_IN_i_31_port, 
      DATA_MEM_IN_i_30_port, DATA_MEM_IN_i_29_port, DATA_MEM_IN_i_28_port, 
      DATA_MEM_IN_i_27_port, DATA_MEM_IN_i_26_port, DATA_MEM_IN_i_25_port, 
      DATA_MEM_IN_i_24_port, DATA_MEM_IN_i_23_port, DATA_MEM_IN_i_22_port, 
      DATA_MEM_IN_i_21_port, DATA_MEM_IN_i_20_port, DATA_MEM_IN_i_19_port, 
      DATA_MEM_IN_i_18_port, DATA_MEM_IN_i_17_port, DATA_MEM_IN_i_16_port, 
      DATA_MEM_IN_i_15_port, DATA_MEM_IN_i_14_port, DATA_MEM_IN_i_13_port, 
      DATA_MEM_IN_i_12_port, DATA_MEM_IN_i_11_port, DATA_MEM_IN_i_10_port, 
      DATA_MEM_IN_i_9_port, DATA_MEM_IN_i_8_port, DATA_MEM_IN_i_7_port, 
      DATA_MEM_IN_i_6_port, DATA_MEM_IN_i_5_port, DATA_MEM_IN_i_4_port, 
      DATA_MEM_IN_i_3_port, DATA_MEM_IN_i_2_port, DATA_MEM_IN_i_1_port, 
      DATA_MEM_IN_i_0_port, dram_data_i_31_port, dram_data_i_30_port, 
      dram_data_i_29_port, dram_data_i_28_port, dram_data_i_27_port, 
      dram_data_i_26_port, dram_data_i_25_port, dram_data_i_24_port, 
      dram_data_i_23_port, dram_data_i_22_port, dram_data_i_21_port, 
      dram_data_i_20_port, dram_data_i_19_port, dram_data_i_18_port, 
      dram_data_i_17_port, dram_data_i_16_port, dram_data_i_15_port, 
      dram_data_i_14_port, dram_data_i_13_port, dram_data_i_12_port, 
      dram_data_i_11_port, dram_data_i_10_port, dram_data_i_9_port, 
      dram_data_i_8_port, dram_data_i_7_port, dram_data_i_6_port, 
      dram_data_i_5_port, dram_data_i_4_port, dram_data_i_3_port, 
      dram_data_i_2_port, dram_data_i_1_port, dram_data_i_0_port, DATA_MEM_WM_i
      , n1, n260, n261, n262, n263, n264, n265, n266, n267, n268, n269, n270, 
      n271, n272, n273, n_2413, n_2414, n_2415, n_2416, n_2417, n_2418, n_2419,
      n_2420, n_2421, n_2422, n_2423, n_2424, n_2425, n_2426, n_2427, n_2428, 
      n_2429, n_2430, n_2431, n_2432, n_2433, n_2434, n_2435, n_2436, n_2437, 
      n_2438, n_2439, n_2440, n_2441, n_2442, n_2443, n_2444, n_2445, n_2446, 
      n_2447, n_2448, n_2449, n_2450, n_2451, n_2452, n_2453, n_2454, n_2455, 
      n_2456, n_2457, n_2458, n_2459, n_2460, n_2461 : std_logic;

begin
   
   DRAM_READNOTWRITE_reg : DFF_X1 port map( D => n270, CK => CLK, Q => 
                           DRAM_READNOTWRITE, QN => n_2413);
   n1 <= '0';
   CU_I : 
                           dlx_cu_MICROCODE_MEM_SIZE62_FUNC_SIZE11_OP_CODE_SIZE6_IR_SIZE32_CW_SIZE15 
                           port map( Clk => CLK, Rst => n271, IR_IN(31) => 
                           IR_31_port, IR_IN(30) => IR_30_port, IR_IN(29) => 
                           IR_29_port, IR_IN(28) => IR_28_port, IR_IN(27) => 
                           IR_27_port, IR_IN(26) => IR_26_port, IR_IN(25) => 
                           IR_25_port, IR_IN(24) => IR_24_port, IR_IN(23) => 
                           IR_23_port, IR_IN(22) => IR_22_port, IR_IN(21) => 
                           IR_21_port, IR_IN(20) => IR_20_port, IR_IN(19) => 
                           IR_19_port, IR_IN(18) => IR_18_port, IR_IN(17) => 
                           IR_17_port, IR_IN(16) => IR_16_port, IR_IN(15) => 
                           IR_15_port, IR_IN(14) => IR_14_port, IR_IN(13) => 
                           IR_13_port, IR_IN(12) => IR_12_port, IR_IN(11) => 
                           IR_11_port, IR_IN(10) => IR_10_port, IR_IN(9) => 
                           IR_9_port, IR_IN(8) => IR_8_port, IR_IN(7) => 
                           IR_7_port, IR_IN(6) => IR_6_port, IR_IN(5) => 
                           IR_5_port, IR_IN(4) => IR_4_port, IR_IN(3) => 
                           IR_3_port, IR_IN(2) => IR_2_port, IR_IN(1) => 
                           IR_1_port, IR_IN(0) => IR_0_port, IR_LATCH_EN => 
                           n_2414, NPC_LATCH_EN => n_2415, RegA_LATCH_EN => 
                           n_2416, RegB_LATCH_EN => n_2417, RegIMM_LATCH_EN => 
                           n_2418, MUXA_SEL => n_2419, MUXB_SEL => n_2420, 
                           ALU_OUTREG_EN => n_2421, EQ_COND => n_2422, 
                           ALU_OPCODE(0) => ALU_OPCODE_i_5_port, ALU_OPCODE(1) 
                           => ALU_OPCODE_i_4_port, ALU_OPCODE(2) => 
                           ALU_OPCODE_i_3_port, ALU_OPCODE(3) => 
                           ALU_OPCODE_i_2_port, ALU_OPCODE(4) => 
                           ALU_OPCODE_i_1_port, ALU_OPCODE(5) => 
                           ALU_OPCODE_i_0_port, signed_unsigned => 
                           signed_unsigned_i, DRAM_WE => n_2423, LMD_LATCH_EN 
                           => n_2424, JUMP_EN => n_2425, PC_LATCH_EN => n_2426,
                           WB_MUX_SEL => n_2427, RF_WE => n_2428, lhi_sel => 
                           lhi_sel_i, sb_op => sb_op_i, s_trap => trap_cs_i, 
                           s_ret => ret_cs_i);
   DTPTH_I : DATAPTH_NBIT32_REG_BIT5 port map( CLK => CLK, RST => n271, PC(31) 
                           => PC_31_port, PC(30) => PC_30_port, PC(29) => 
                           PC_29_port, PC(28) => PC_28_port, PC(27) => 
                           PC_27_port, PC(26) => PC_26_port, PC(25) => 
                           PC_25_port, PC(24) => PC_24_port, PC(23) => 
                           PC_23_port, PC(22) => PC_22_port, PC(21) => 
                           PC_21_port, PC(20) => PC_20_port, PC(19) => 
                           PC_19_port, PC(18) => PC_18_port, PC(17) => 
                           PC_17_port, PC(16) => PC_16_port, PC(15) => 
                           PC_15_port, PC(14) => PC_14_port, PC(13) => 
                           PC_13_port, PC(12) => PC_12_port, PC(11) => 
                           PC_11_port, PC(10) => PC_10_port, PC(9) => PC_9_port
                           , PC(8) => PC_8_port, PC(7) => PC_7_port, PC(6) => 
                           PC_6_port, PC(5) => PC_5_port, PC(4) => PC_4_port, 
                           PC(3) => PC_3_port, PC(2) => PC_2_port, PC(1) => 
                           PC_1_port, PC(0) => PC_0_port, IR(31) => IR_31_port,
                           IR(30) => IR_30_port, IR(29) => IR_29_port, IR(28) 
                           => IR_28_port, IR(27) => IR_27_port, IR(26) => 
                           IR_26_port, IR(25) => IR_25_port, IR(24) => 
                           IR_24_port, IR(23) => IR_23_port, IR(22) => 
                           IR_22_port, IR(21) => IR_21_port, IR(20) => 
                           IR_20_port, IR(19) => IR_19_port, IR(18) => 
                           IR_18_port, IR(17) => IR_17_port, IR(16) => 
                           IR_16_port, IR(15) => IR_15_port, IR(14) => 
                           IR_14_port, IR(13) => IR_13_port, IR(12) => 
                           IR_12_port, IR(11) => IR_11_port, IR(10) => 
                           IR_10_port, IR(9) => IR_9_port, IR(8) => IR_8_port, 
                           IR(7) => IR_7_port, IR(6) => IR_6_port, IR(5) => 
                           IR_5_port, IR(4) => IR_4_port, IR(3) => IR_3_port, 
                           IR(2) => IR_2_port, IR(1) => IR_1_port, IR(0) => 
                           IR_0_port, PC_OUT(31) => n_2429, PC_OUT(30) => 
                           n_2430, PC_OUT(29) => n_2431, PC_OUT(28) => n_2432, 
                           PC_OUT(27) => n_2433, PC_OUT(26) => n_2434, 
                           PC_OUT(25) => n_2435, PC_OUT(24) => n_2436, 
                           PC_OUT(23) => n_2437, PC_OUT(22) => n_2438, 
                           PC_OUT(21) => n_2439, PC_OUT(20) => n_2440, 
                           PC_OUT(19) => n_2441, PC_OUT(18) => n_2442, 
                           PC_OUT(17) => n_2443, PC_OUT(16) => n_2444, 
                           PC_OUT(15) => n_2445, PC_OUT(14) => n_2446, 
                           PC_OUT(13) => n_2447, PC_OUT(12) => n_2448, 
                           PC_OUT(11) => n_2449, PC_OUT(10) => n_2450, 
                           PC_OUT(9) => n_2451, PC_OUT(8) => n_2452, PC_OUT(7) 
                           => n_2453, PC_OUT(6) => n_2454, PC_OUT(5) => n_2455,
                           PC_OUT(4) => n_2456, PC_OUT(3) => n_2457, PC_OUT(2) 
                           => n_2458, PC_OUT(1) => n_2459, PC_OUT(0) => n_2460,
                           NPC_LATCH_EN => NPC_LATCH_EN_i, ir_LATCH_EN => 
                           IR_LATCH_EN_i, signed_op => signed_unsigned_i, 
                           trap_cs => trap_cs_i, ret_cs => ret_cs_i, RF1 => 
                           RegA_LATCH_EN_i, RF2 => RegB_LATCH_EN_i, WF1 => 
                           RF_WE_i, regImm_LATCH_EN => RegIMM_LATCH_EN_i, S1 =>
                           MUXA_SEL_i, S2 => MUXB_SEL_i, EN2 => ALU_OUTREG_EN_i
                           , lhi_sel => lhi_sel_i, jump_en => JUMP_EN_i, 
                           branch_cond => EQ_COND_i, sb_op => sb_op_i, RM => 
                           LMD_LATCH_EN_i, WM => DRAM_WE_i, EN3 => 
                           PC_LATCH_EN_i, S3 => WB_MUX_SEL_i, 
                           instruction_alu(0) => ALU_OPCODE_i_5_port, 
                           instruction_alu(1) => ALU_OPCODE_i_4_port, 
                           instruction_alu(2) => ALU_OPCODE_i_3_port, 
                           instruction_alu(3) => ALU_OPCODE_i_2_port, 
                           instruction_alu(4) => ALU_OPCODE_i_1_port, 
                           instruction_alu(5) => ALU_OPCODE_i_0_port, 
                           DATA_MEM_ADDR(31) => DRAM_ADDRESS(31), 
                           DATA_MEM_ADDR(30) => DRAM_ADDRESS(30), 
                           DATA_MEM_ADDR(29) => DRAM_ADDRESS(29), 
                           DATA_MEM_ADDR(28) => DRAM_ADDRESS(28), 
                           DATA_MEM_ADDR(27) => DRAM_ADDRESS(27), 
                           DATA_MEM_ADDR(26) => DRAM_ADDRESS(26), 
                           DATA_MEM_ADDR(25) => DRAM_ADDRESS(25), 
                           DATA_MEM_ADDR(24) => DRAM_ADDRESS(24), 
                           DATA_MEM_ADDR(23) => DRAM_ADDRESS(23), 
                           DATA_MEM_ADDR(22) => DRAM_ADDRESS(22), 
                           DATA_MEM_ADDR(21) => DRAM_ADDRESS(21), 
                           DATA_MEM_ADDR(20) => DRAM_ADDRESS(20), 
                           DATA_MEM_ADDR(19) => DRAM_ADDRESS(19), 
                           DATA_MEM_ADDR(18) => DRAM_ADDRESS(18), 
                           DATA_MEM_ADDR(17) => DRAM_ADDRESS(17), 
                           DATA_MEM_ADDR(16) => DRAM_ADDRESS(16), 
                           DATA_MEM_ADDR(15) => DRAM_ADDRESS(15), 
                           DATA_MEM_ADDR(14) => DRAM_ADDRESS(14), 
                           DATA_MEM_ADDR(13) => DRAM_ADDRESS(13), 
                           DATA_MEM_ADDR(12) => DRAM_ADDRESS(12), 
                           DATA_MEM_ADDR(11) => DRAM_ADDRESS(11), 
                           DATA_MEM_ADDR(10) => DRAM_ADDRESS(10), 
                           DATA_MEM_ADDR(9) => DRAM_ADDRESS(9), 
                           DATA_MEM_ADDR(8) => DRAM_ADDRESS(8), 
                           DATA_MEM_ADDR(7) => DRAM_ADDRESS(7), 
                           DATA_MEM_ADDR(6) => DRAM_ADDRESS(6), 
                           DATA_MEM_ADDR(5) => DRAM_ADDRESS(5), 
                           DATA_MEM_ADDR(4) => DRAM_ADDRESS(4), 
                           DATA_MEM_ADDR(3) => DRAM_ADDRESS(3), 
                           DATA_MEM_ADDR(2) => DRAM_ADDRESS(2), 
                           DATA_MEM_ADDR(1) => DRAM_ADDRESS(1), 
                           DATA_MEM_ADDR(0) => DRAM_ADDRESS(0), DATA_MEM_IN(31)
                           => DATA_MEM_IN_i_31_port, DATA_MEM_IN(30) => 
                           DATA_MEM_IN_i_30_port, DATA_MEM_IN(29) => 
                           DATA_MEM_IN_i_29_port, DATA_MEM_IN(28) => 
                           DATA_MEM_IN_i_28_port, DATA_MEM_IN(27) => 
                           DATA_MEM_IN_i_27_port, DATA_MEM_IN(26) => 
                           DATA_MEM_IN_i_26_port, DATA_MEM_IN(25) => 
                           DATA_MEM_IN_i_25_port, DATA_MEM_IN(24) => 
                           DATA_MEM_IN_i_24_port, DATA_MEM_IN(23) => 
                           DATA_MEM_IN_i_23_port, DATA_MEM_IN(22) => 
                           DATA_MEM_IN_i_22_port, DATA_MEM_IN(21) => 
                           DATA_MEM_IN_i_21_port, DATA_MEM_IN(20) => 
                           DATA_MEM_IN_i_20_port, DATA_MEM_IN(19) => 
                           DATA_MEM_IN_i_19_port, DATA_MEM_IN(18) => 
                           DATA_MEM_IN_i_18_port, DATA_MEM_IN(17) => 
                           DATA_MEM_IN_i_17_port, DATA_MEM_IN(16) => 
                           DATA_MEM_IN_i_16_port, DATA_MEM_IN(15) => 
                           DATA_MEM_IN_i_15_port, DATA_MEM_IN(14) => 
                           DATA_MEM_IN_i_14_port, DATA_MEM_IN(13) => 
                           DATA_MEM_IN_i_13_port, DATA_MEM_IN(12) => 
                           DATA_MEM_IN_i_12_port, DATA_MEM_IN(11) => 
                           DATA_MEM_IN_i_11_port, DATA_MEM_IN(10) => 
                           DATA_MEM_IN_i_10_port, DATA_MEM_IN(9) => 
                           DATA_MEM_IN_i_9_port, DATA_MEM_IN(8) => 
                           DATA_MEM_IN_i_8_port, DATA_MEM_IN(7) => 
                           DATA_MEM_IN_i_7_port, DATA_MEM_IN(6) => 
                           DATA_MEM_IN_i_6_port, DATA_MEM_IN(5) => 
                           DATA_MEM_IN_i_5_port, DATA_MEM_IN(4) => 
                           DATA_MEM_IN_i_4_port, DATA_MEM_IN(3) => 
                           DATA_MEM_IN_i_3_port, DATA_MEM_IN(2) => 
                           DATA_MEM_IN_i_2_port, DATA_MEM_IN(1) => 
                           DATA_MEM_IN_i_1_port, DATA_MEM_IN(0) => 
                           DATA_MEM_IN_i_0_port, DATA_MEM_OUT(31) => 
                           dram_data_i_31_port, DATA_MEM_OUT(30) => 
                           dram_data_i_30_port, DATA_MEM_OUT(29) => 
                           dram_data_i_29_port, DATA_MEM_OUT(28) => 
                           dram_data_i_28_port, DATA_MEM_OUT(27) => 
                           dram_data_i_27_port, DATA_MEM_OUT(26) => 
                           dram_data_i_26_port, DATA_MEM_OUT(25) => 
                           dram_data_i_25_port, DATA_MEM_OUT(24) => 
                           dram_data_i_24_port, DATA_MEM_OUT(23) => 
                           dram_data_i_23_port, DATA_MEM_OUT(22) => 
                           dram_data_i_22_port, DATA_MEM_OUT(21) => 
                           dram_data_i_21_port, DATA_MEM_OUT(20) => 
                           dram_data_i_20_port, DATA_MEM_OUT(19) => 
                           dram_data_i_19_port, DATA_MEM_OUT(18) => 
                           dram_data_i_18_port, DATA_MEM_OUT(17) => 
                           dram_data_i_17_port, DATA_MEM_OUT(16) => 
                           dram_data_i_16_port, DATA_MEM_OUT(15) => 
                           dram_data_i_15_port, DATA_MEM_OUT(14) => 
                           dram_data_i_14_port, DATA_MEM_OUT(13) => 
                           dram_data_i_13_port, DATA_MEM_OUT(12) => 
                           dram_data_i_12_port, DATA_MEM_OUT(11) => 
                           dram_data_i_11_port, DATA_MEM_OUT(10) => 
                           dram_data_i_10_port, DATA_MEM_OUT(9) => 
                           dram_data_i_9_port, DATA_MEM_OUT(8) => 
                           dram_data_i_8_port, DATA_MEM_OUT(7) => 
                           dram_data_i_7_port, DATA_MEM_OUT(6) => 
                           dram_data_i_6_port, DATA_MEM_OUT(5) => 
                           dram_data_i_5_port, DATA_MEM_OUT(4) => 
                           dram_data_i_4_port, DATA_MEM_OUT(3) => 
                           dram_data_i_3_port, DATA_MEM_OUT(2) => 
                           dram_data_i_2_port, DATA_MEM_OUT(1) => 
                           dram_data_i_1_port, DATA_MEM_OUT(0) => 
                           dram_data_i_0_port, DATA_MEM_ENABLE => DRAM_ISSUE, 
                           DATA_MEM_RM => n_2461, DATA_MEM_WM => DATA_MEM_WM_i)
                           ;
   DRAM_DATA_tri_32_inst : TBUF_X1 port map( A => n1, EN => n266, Z => 
                           DRAM_DATA(32));
   DRAM_DATA_tri_33_inst : TBUF_X1 port map( A => n1, EN => n264, Z => 
                           DRAM_DATA(33));
   DRAM_DATA_tri_34_inst : TBUF_X1 port map( A => n1, EN => n266, Z => 
                           DRAM_DATA(34));
   DRAM_DATA_tri_35_inst : TBUF_X1 port map( A => n1, EN => n264, Z => 
                           DRAM_DATA(35));
   DRAM_DATA_tri_36_inst : TBUF_X1 port map( A => n1, EN => n266, Z => 
                           DRAM_DATA(36));
   DRAM_DATA_tri_37_inst : TBUF_X1 port map( A => n1, EN => n264, Z => 
                           DRAM_DATA(37));
   DRAM_DATA_tri_38_inst : TBUF_X1 port map( A => n1, EN => n266, Z => 
                           DRAM_DATA(38));
   DRAM_DATA_tri_39_inst : TBUF_X1 port map( A => n1, EN => n264, Z => 
                           DRAM_DATA(39));
   DRAM_DATA_tri_40_inst : TBUF_X1 port map( A => n1, EN => n264, Z => 
                           DRAM_DATA(40));
   DRAM_DATA_tri_41_inst : TBUF_X1 port map( A => n1, EN => n267, Z => 
                           DRAM_DATA(41));
   DRAM_DATA_tri_42_inst : TBUF_X1 port map( A => n1, EN => n264, Z => 
                           DRAM_DATA(42));
   DRAM_DATA_tri_43_inst : TBUF_X1 port map( A => n1, EN => n267, Z => 
                           DRAM_DATA(43));
   DRAM_DATA_tri_44_inst : TBUF_X1 port map( A => n1, EN => n264, Z => 
                           DRAM_DATA(44));
   DRAM_DATA_tri_45_inst : TBUF_X1 port map( A => n1, EN => n267, Z => 
                           DRAM_DATA(45));
   DRAM_DATA_tri_46_inst : TBUF_X1 port map( A => n1, EN => n263, Z => 
                           DRAM_DATA(46));
   DRAM_DATA_tri_47_inst : TBUF_X1 port map( A => n1, EN => n267, Z => 
                           DRAM_DATA(47));
   DRAM_DATA_tri_48_inst : TBUF_X1 port map( A => n1, EN => n263, Z => 
                           DRAM_DATA(48));
   DRAM_DATA_tri_49_inst : TBUF_X1 port map( A => n1, EN => n267, Z => 
                           DRAM_DATA(49));
   DRAM_DATA_tri_50_inst : TBUF_X1 port map( A => n1, EN => n267, Z => 
                           DRAM_DATA(50));
   DRAM_DATA_tri_51_inst : TBUF_X1 port map( A => n1, EN => n263, Z => 
                           DRAM_DATA(51));
   DRAM_DATA_tri_52_inst : TBUF_X1 port map( A => n1, EN => n267, Z => 
                           DRAM_DATA(52));
   DRAM_DATA_tri_53_inst : TBUF_X1 port map( A => n1, EN => n263, Z => 
                           DRAM_DATA(53));
   DRAM_DATA_tri_54_inst : TBUF_X1 port map( A => n1, EN => n267, Z => 
                           DRAM_DATA(54));
   DRAM_DATA_tri_55_inst : TBUF_X1 port map( A => n1, EN => n263, Z => 
                           DRAM_DATA(55));
   DRAM_DATA_tri_56_inst : TBUF_X1 port map( A => n1, EN => n267, Z => 
                           DRAM_DATA(56));
   DRAM_DATA_tri_57_inst : TBUF_X1 port map( A => n1, EN => n263, Z => 
                           DRAM_DATA(57));
   DRAM_DATA_tri_58_inst : TBUF_X1 port map( A => n1, EN => n267, Z => 
                           DRAM_DATA(58));
   DRAM_DATA_tri_59_inst : TBUF_X1 port map( A => n1, EN => n263, Z => 
                           DRAM_DATA(59));
   DRAM_DATA_tri_60_inst : TBUF_X1 port map( A => n1, EN => n263, Z => 
                           DRAM_DATA(60));
   DRAM_DATA_tri_61_inst : TBUF_X1 port map( A => n1, EN => n268, Z => 
                           DRAM_DATA(61));
   DRAM_DATA_tri_62_inst : TBUF_X1 port map( A => n1, EN => n263, Z => 
                           DRAM_DATA(62));
   DRAM_DATA_tri_63_inst : TBUF_X1 port map( A => n1, EN => n268, Z => 
                           DRAM_DATA(63));
   DRAM_DATA_tri_0_inst : TBUF_X1 port map( A => DATA_MEM_IN_i_0_port, EN => 
                           n265, Z => DRAM_DATA(0));
   DRAM_DATA_tri_1_inst : TBUF_X1 port map( A => DATA_MEM_IN_i_1_port, EN => 
                           n266, Z => DRAM_DATA(1));
   DRAM_DATA_tri_2_inst : TBUF_X1 port map( A => DATA_MEM_IN_i_2_port, EN => 
                           n264, Z => DRAM_DATA(2));
   DRAM_DATA_tri_3_inst : TBUF_X1 port map( A => DATA_MEM_IN_i_3_port, EN => 
                           n267, Z => DRAM_DATA(3));
   DRAM_DATA_tri_4_inst : TBUF_X1 port map( A => DATA_MEM_IN_i_4_port, EN => 
                           n263, Z => DRAM_DATA(4));
   DRAM_DATA_tri_5_inst : TBUF_X1 port map( A => DATA_MEM_IN_i_5_port, EN => 
                           n267, Z => DRAM_DATA(5));
   DRAM_DATA_tri_6_inst : TBUF_X1 port map( A => DATA_MEM_IN_i_6_port, EN => 
                           n263, Z => DRAM_DATA(6));
   DRAM_DATA_tri_7_inst : TBUF_X1 port map( A => DATA_MEM_IN_i_7_port, EN => 
                           n268, Z => DRAM_DATA(7));
   DRAM_DATA_tri_8_inst : TBUF_X1 port map( A => DATA_MEM_IN_i_8_port, EN => 
                           n263, Z => DRAM_DATA(8));
   DRAM_DATA_tri_9_inst : TBUF_X1 port map( A => DATA_MEM_IN_i_9_port, EN => 
                           n268, Z => DRAM_DATA(9));
   DRAM_DATA_tri_10_inst : TBUF_X1 port map( A => DATA_MEM_IN_i_10_port, EN => 
                           n265, Z => DRAM_DATA(10));
   DRAM_DATA_tri_11_inst : TBUF_X1 port map( A => DATA_MEM_IN_i_11_port, EN => 
                           n265, Z => DRAM_DATA(11));
   DRAM_DATA_tri_12_inst : TBUF_X1 port map( A => DATA_MEM_IN_i_12_port, EN => 
                           n265, Z => DRAM_DATA(12));
   DRAM_DATA_tri_13_inst : TBUF_X1 port map( A => DATA_MEM_IN_i_13_port, EN => 
                           n265, Z => DRAM_DATA(13));
   DRAM_DATA_tri_14_inst : TBUF_X1 port map( A => DATA_MEM_IN_i_14_port, EN => 
                           n265, Z => DRAM_DATA(14));
   DRAM_DATA_tri_15_inst : TBUF_X1 port map( A => DATA_MEM_IN_i_15_port, EN => 
                           n265, Z => DRAM_DATA(15));
   DRAM_DATA_tri_16_inst : TBUF_X1 port map( A => DATA_MEM_IN_i_16_port, EN => 
                           n265, Z => DRAM_DATA(16));
   DRAM_DATA_tri_17_inst : TBUF_X1 port map( A => DATA_MEM_IN_i_17_port, EN => 
                           n265, Z => DRAM_DATA(17));
   DRAM_DATA_tri_18_inst : TBUF_X1 port map( A => DATA_MEM_IN_i_18_port, EN => 
                           n266, Z => DRAM_DATA(18));
   DRAM_DATA_tri_19_inst : TBUF_X1 port map( A => DATA_MEM_IN_i_19_port, EN => 
                           n265, Z => DRAM_DATA(19));
   DRAM_DATA_tri_20_inst : TBUF_X1 port map( A => DATA_MEM_IN_i_20_port, EN => 
                           n265, Z => DRAM_DATA(20));
   DRAM_DATA_tri_21_inst : TBUF_X1 port map( A => DATA_MEM_IN_i_21_port, EN => 
                           n266, Z => DRAM_DATA(21));
   DRAM_DATA_tri_22_inst : TBUF_X1 port map( A => DATA_MEM_IN_i_22_port, EN => 
                           n265, Z => DRAM_DATA(22));
   DRAM_DATA_tri_23_inst : TBUF_X1 port map( A => DATA_MEM_IN_i_23_port, EN => 
                           n266, Z => DRAM_DATA(23));
   DRAM_DATA_tri_24_inst : TBUF_X1 port map( A => DATA_MEM_IN_i_24_port, EN => 
                           n264, Z => DRAM_DATA(24));
   DRAM_DATA_tri_25_inst : TBUF_X1 port map( A => DATA_MEM_IN_i_25_port, EN => 
                           n266, Z => DRAM_DATA(25));
   DRAM_DATA_tri_26_inst : TBUF_X1 port map( A => DATA_MEM_IN_i_26_port, EN => 
                           n264, Z => DRAM_DATA(26));
   DRAM_DATA_tri_27_inst : TBUF_X1 port map( A => DATA_MEM_IN_i_27_port, EN => 
                           n266, Z => DRAM_DATA(27));
   DRAM_DATA_tri_28_inst : TBUF_X1 port map( A => DATA_MEM_IN_i_28_port, EN => 
                           n264, Z => DRAM_DATA(28));
   DRAM_DATA_tri_29_inst : TBUF_X1 port map( A => DATA_MEM_IN_i_29_port, EN => 
                           n266, Z => DRAM_DATA(29));
   DRAM_DATA_tri_30_inst : TBUF_X1 port map( A => DATA_MEM_IN_i_30_port, EN => 
                           n266, Z => DRAM_DATA(30));
   DRAM_DATA_tri_31_inst : TBUF_X1 port map( A => DATA_MEM_IN_i_31_port, EN => 
                           n264, Z => DRAM_DATA(31));
   U198 : BUF_X1 port map( A => n260, Z => n263);
   U199 : BUF_X1 port map( A => n261, Z => n267);
   U200 : BUF_X1 port map( A => n260, Z => n264);
   U201 : BUF_X1 port map( A => n261, Z => n266);
   U202 : BUF_X1 port map( A => n260, Z => n265);
   U203 : BUF_X1 port map( A => n261, Z => n268);
   U204 : BUF_X1 port map( A => n262, Z => n269);
   U205 : AND2_X1 port map( A1 => DRAM_DATA(63), A2 => n269, ZN => 
                           dram_data_i_31_port);
   U206 : AND2_X1 port map( A1 => DRAM_DATA(40), A2 => n270, ZN => 
                           dram_data_i_8_port);
   U207 : AND2_X1 port map( A1 => DRAM_DATA(41), A2 => n270, ZN => 
                           dram_data_i_9_port);
   U208 : AND2_X1 port map( A1 => DRAM_DATA(42), A2 => n268, ZN => 
                           dram_data_i_10_port);
   U209 : AND2_X1 port map( A1 => DRAM_DATA(43), A2 => n268, ZN => 
                           dram_data_i_11_port);
   U210 : AND2_X1 port map( A1 => DRAM_DATA(44), A2 => n268, ZN => 
                           dram_data_i_12_port);
   U211 : AND2_X1 port map( A1 => DRAM_DATA(45), A2 => n268, ZN => 
                           dram_data_i_13_port);
   U212 : AND2_X1 port map( A1 => DRAM_DATA(46), A2 => n268, ZN => 
                           dram_data_i_14_port);
   U213 : AND2_X1 port map( A1 => DRAM_DATA(47), A2 => n268, ZN => 
                           dram_data_i_15_port);
   U214 : AND2_X1 port map( A1 => DRAM_DATA(52), A2 => n269, ZN => 
                           dram_data_i_20_port);
   U215 : AND2_X1 port map( A1 => DRAM_DATA(53), A2 => n269, ZN => 
                           dram_data_i_21_port);
   U216 : AND2_X1 port map( A1 => DRAM_DATA(54), A2 => n269, ZN => 
                           dram_data_i_22_port);
   U217 : AND2_X1 port map( A1 => DRAM_DATA(55), A2 => n269, ZN => 
                           dram_data_i_23_port);
   U218 : AND2_X1 port map( A1 => DRAM_DATA(56), A2 => n269, ZN => 
                           dram_data_i_24_port);
   U219 : AND2_X1 port map( A1 => DRAM_DATA(57), A2 => n269, ZN => 
                           dram_data_i_25_port);
   U220 : AND2_X1 port map( A1 => DRAM_DATA(58), A2 => n269, ZN => 
                           dram_data_i_26_port);
   U221 : AND2_X1 port map( A1 => DRAM_DATA(59), A2 => n269, ZN => 
                           dram_data_i_27_port);
   U222 : AND2_X1 port map( A1 => DRAM_DATA(60), A2 => n269, ZN => 
                           dram_data_i_28_port);
   U223 : AND2_X1 port map( A1 => DRAM_DATA(61), A2 => n269, ZN => 
                           dram_data_i_29_port);
   U224 : AND2_X1 port map( A1 => DRAM_DATA(62), A2 => n269, ZN => 
                           dram_data_i_30_port);
   U225 : AND2_X1 port map( A1 => DRAM_DATA(48), A2 => n268, ZN => 
                           dram_data_i_16_port);
   U226 : AND2_X1 port map( A1 => DRAM_DATA(49), A2 => n268, ZN => 
                           dram_data_i_17_port);
   U227 : AND2_X1 port map( A1 => DRAM_DATA(50), A2 => n268, ZN => 
                           dram_data_i_18_port);
   U228 : AND2_X1 port map( A1 => DRAM_DATA(51), A2 => n269, ZN => 
                           dram_data_i_19_port);
   U229 : BUF_X1 port map( A => n272, Z => n271);
   U230 : BUF_X1 port map( A => RST, Z => n272);
   U231 : AND2_X1 port map( A1 => DRAM_DATA(32), A2 => n268, ZN => 
                           dram_data_i_0_port);
   U232 : AND2_X1 port map( A1 => DRAM_DATA(33), A2 => n268, ZN => 
                           dram_data_i_1_port);
   U233 : AND2_X1 port map( A1 => DRAM_DATA(34), A2 => n269, ZN => 
                           dram_data_i_2_port);
   U234 : AND2_X1 port map( A1 => DRAM_DATA(35), A2 => n269, ZN => 
                           dram_data_i_3_port);
   U235 : AND2_X1 port map( A1 => DRAM_DATA(36), A2 => n270, ZN => 
                           dram_data_i_4_port);
   U236 : AND2_X1 port map( A1 => DRAM_DATA(37), A2 => n269, ZN => 
                           dram_data_i_5_port);
   U237 : AND2_X1 port map( A1 => DRAM_DATA(38), A2 => n270, ZN => 
                           dram_data_i_6_port);
   U238 : AND2_X1 port map( A1 => DRAM_DATA(39), A2 => n270, ZN => 
                           dram_data_i_7_port);
   U239 : INV_X1 port map( A => DATA_MEM_WM_i, ZN => n273);
   IR_0_port <= '0';
   IR_1_port <= '0';
   IR_2_port <= '0';
   IR_3_port <= '0';
   IR_4_port <= '0';
   IR_5_port <= '0';
   IR_6_port <= '0';
   IR_7_port <= '0';
   IR_8_port <= '0';
   IR_9_port <= '0';
   IR_10_port <= '0';
   IR_11_port <= '0';
   IR_12_port <= '0';
   IR_13_port <= '0';
   IR_14_port <= '0';
   IR_15_port <= '0';
   IR_16_port <= '0';
   IR_17_port <= '0';
   IR_18_port <= '0';
   IR_19_port <= '0';
   IR_20_port <= '0';
   IR_21_port <= '0';
   IR_22_port <= '0';
   IR_23_port <= '0';
   IR_24_port <= '0';
   IR_25_port <= '0';
   IR_26_port <= '0';
   IR_27_port <= '0';
   IR_28_port <= '0';
   IR_29_port <= '0';
   IR_30_port <= '0';
   IR_31_port <= '0';
   PC_0_port <= '0';
   IRAM_ADDRESS(0) <= '0';
   PC_1_port <= '0';
   IRAM_ADDRESS(1) <= '0';
   PC_2_port <= '0';
   IRAM_ADDRESS(2) <= '0';
   PC_3_port <= '0';
   IRAM_ADDRESS(3) <= '0';
   PC_4_port <= '0';
   IRAM_ADDRESS(4) <= '0';
   PC_5_port <= '0';
   IRAM_ADDRESS(5) <= '0';
   PC_6_port <= '0';
   IRAM_ADDRESS(6) <= '0';
   PC_7_port <= '0';
   IRAM_ADDRESS(7) <= '0';
   PC_8_port <= '0';
   IRAM_ADDRESS(8) <= '0';
   PC_9_port <= '0';
   IRAM_ADDRESS(9) <= '0';
   PC_10_port <= '0';
   IRAM_ADDRESS(10) <= '0';
   PC_11_port <= '0';
   IRAM_ADDRESS(11) <= '0';
   PC_12_port <= '0';
   IRAM_ADDRESS(12) <= '0';
   PC_13_port <= '0';
   IRAM_ADDRESS(13) <= '0';
   PC_14_port <= '0';
   IRAM_ADDRESS(14) <= '0';
   PC_15_port <= '0';
   IRAM_ADDRESS(15) <= '0';
   PC_16_port <= '0';
   IRAM_ADDRESS(16) <= '0';
   PC_17_port <= '0';
   IRAM_ADDRESS(17) <= '0';
   PC_18_port <= '0';
   IRAM_ADDRESS(18) <= '0';
   PC_19_port <= '0';
   IRAM_ADDRESS(19) <= '0';
   PC_20_port <= '0';
   IRAM_ADDRESS(20) <= '0';
   PC_21_port <= '0';
   IRAM_ADDRESS(21) <= '0';
   PC_22_port <= '0';
   IRAM_ADDRESS(22) <= '0';
   PC_23_port <= '0';
   IRAM_ADDRESS(23) <= '0';
   PC_24_port <= '0';
   IRAM_ADDRESS(24) <= '0';
   PC_25_port <= '0';
   IRAM_ADDRESS(25) <= '0';
   PC_26_port <= '0';
   IRAM_ADDRESS(26) <= '0';
   PC_27_port <= '0';
   IRAM_ADDRESS(27) <= '0';
   PC_28_port <= '0';
   IRAM_ADDRESS(28) <= '0';
   PC_29_port <= '0';
   IRAM_ADDRESS(29) <= '0';
   PC_30_port <= '0';
   IRAM_ADDRESS(30) <= '0';
   PC_31_port <= '0';
   IRAM_ADDRESS(31) <= '0';
   U336 : CLKBUF_X1 port map( A => n273, Z => n260);
   U337 : CLKBUF_X1 port map( A => n273, Z => n261);
   U338 : CLKBUF_X1 port map( A => n273, Z => n262);
   U339 : CLKBUF_X1 port map( A => n262, Z => n270);
   RF_WE_i <= '0';
   WB_MUX_SEL_i <= '0';
   PC_LATCH_EN_i <= '0';
   JUMP_EN_i <= '0';
   LMD_LATCH_EN_i <= '0';
   DRAM_WE_i <= '0';
   EQ_COND_i <= '0';
   ALU_OUTREG_EN_i <= '0';
   MUXB_SEL_i <= '0';
   MUXA_SEL_i <= '0';
   RegIMM_LATCH_EN_i <= '0';
   RegB_LATCH_EN_i <= '0';
   RegA_LATCH_EN_i <= '0';
   NPC_LATCH_EN_i <= '0';
   IR_LATCH_EN_i <= '0';

end SYN_dlx_rtl;
